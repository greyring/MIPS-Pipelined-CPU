`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    00:15:45 12/12/2017 
// Design Name: 
// Module Name:    tlb_mem 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module tlb_mem(
	input clk,
	input rst
	
	
	
    );
parameter DATA_SIZE = 1;


endmodule
