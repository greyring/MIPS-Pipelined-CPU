//	`define DEBUG