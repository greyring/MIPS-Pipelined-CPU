`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    19:28:31 09/04/2017 
// Design Name: 
// Module Name:    top 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
`include "define.vh"
module top(
	input clk200P,
	input clk200N,
	`ifdef DEBUG
	input clk_100mhz,
	input clk_uart,
	input [4:0]int_,
	`endif
	
    output [4:0] btn_x,
	 input [4:0] btn_y,
	 input [15:0] switch,
    input RSTN,
    
   output led_clk,
   output led_do,
   output led_pen,
   output seg_clk,
   output seg_do,
   output seg_pen,
	
	output [3:0]vga_red,
	output [3:0]vga_green,
	output [3:0]vga_blue,
	output vga_h_sync,
	output vga_v_sync,
	
	input ps2_clk,
	input ps2_dat,
	
	input uart_rx,
	output uart_tx
    );
`ifdef DEBUG
reg [31:0]Div = 32'b0;
always @(posedge clk_100mhz)
	Div <= Div+1;
`else
wire clk_100mhz;
wire [31:0]Div;
clk_gen_sword clk_gen(
    .clk_pad_p(clk200P), 
    .clk_pad_n(clk200N), 
    .clk_100m(clk_100mhz), 
    .clk_50m(), 
    .clk_25m(), 
    .clk_10m(), 
    .Div(Div), 
    .locked()
    );
`endif

wire [15:0]SW_OK;
wire [24:0]BTN_OK;
wire rst;
input_switch_btn Input_switch_btn(
    .clk(clk_100mhz), 
    .RSTN(RSTN), 
    .switch(switch), 
    .btn_x(btn_x), 
    .btn_y(btn_y), 
    .sw_ok(SW_OK), 
    .btn_ok(BTN_OK),
	 .cr(),
	 .rst(rst)
    );

wire Clk_CPU;
assign Clk_CPU = SW_OK[2]? Div[24]:Div[0];//50m�е�죿

wire [31:0]addr_bus;
wire [31:0]data_bus;
wire [5:0]ctrl_bus;
wire  en_TEXTS, en_DATAS, en_BIOS, en_vga_reg, en_cursor_reg, en_textRAM, 
		en_graphRAM, en_DRAM, en_SEG, en_keyboard, en_switch, en_led, en_dma, en_dmaRAM, en_others;//en_SRAM,
addr_decoder Addr_decoder(
    .addr(addr_bus), 
    .en_TEXTS(en_TEXTS), .en_DATAS(en_DATAS), .en_BIOS(en_BIOS), .en_vga_reg(en_vga_reg),     
	 .en_cursor_reg(en_cursor_reg), .en_textRAM(en_textRAM),     
	 .en_graphRAM(en_graphRAM), .en_DRAM(en_DRAM), .en_SEG(en_SEG), 
	 .en_keyboard(en_keyboard), .en_switch(en_switch), .en_led(en_led),
	 .en_dma(en_dma), .en_dmaRAM(en_dmaRAM),
    .en_others(en_others)
    );//.en_SRAM(en_SRAM),
/*
wire [31:0]SRAM_addr, SRAM_wdata, SRAM_rdata;
wire SRAM_r;
wire [3:0]SRAM_w;
bus_interface SRAM(
    .enable(en_SRAM), 
    .addr(addr_bus), .data(data_bus), .r(ctrl_bus[0]), .w(ctrl_bus[4:1]), .ready(ctrl_bus[5]), 
    .addr_(SRAM_addr), .wdata(SRAM_wdata), .rdata(SRAM_rdata), 
	 .r_(SRAM_r), .w_(SRAM_w), .ready_(1'b1)
    );
*/
wire [31:0]TEXTS_baddr, TEXTS_bwdata, TEXTS_brdata;
wire TEXTS_br;
wire [3:0]TEXTS_bw;
bus_interface TEXTS(
    .enable(en_TEXTS), 
    .addr(addr_bus), .data(data_bus), .r(ctrl_bus[0]), .w(ctrl_bus[4:1]), .ready(ctrl_bus[5]), 
    .addr_(TEXTS_baddr), .wdata(TEXTS_bwdata), .rdata(TEXTS_brdata), 
	 .r_(TEXTS_br), .w_(TEXTS_bw), .ready_(1'b1)
    );
wire [31:0]DATAS_baddr, DATAS_bwdata, DATAS_brdata;
wire DATAS_br;
wire [3:0]DATAS_bw;
bus_interface DATAS(
    .enable(en_DATAS), 
    .addr(addr_bus), .data(data_bus), .r(ctrl_bus[0]), .w(ctrl_bus[4:1]), .ready(ctrl_bus[5]), 
    .addr_(DATAS_baddr), .wdata(DATAS_bwdata), .rdata(DATAS_brdata), 
	 .r_(DATAS_br), .w_(DATAS_bw), .ready_(1'b1)
    );
wire [31:0]vga_reg_wdata, vga_reg_rdata;
wire vga_reg_r;
wire [3:0]vga_reg_w;
bus_interface VGA_REG(
    .enable(en_vga_reg), 
    .addr(addr_bus), .data(data_bus), .r(ctrl_bus[0]), .w(ctrl_bus[4:1]), .ready(ctrl_bus[5]), 
    .addr_(), .wdata(vga_reg_wdata), .rdata(vga_reg_rdata), 
	 .r_(vga_reg_r), .w_(vga_reg_w), .ready_(1'b1)
    );
wire [31:0]vga_cursor_wdata, vga_cursor_rdata;
wire vga_cursor_r;
wire [3:0]vga_cursor_w;
bus_interface VGA_CURSOR(
    .enable(en_cursor_reg), 
    .addr(addr_bus), .data(data_bus), .r(ctrl_bus[0]), .w(ctrl_bus[4:1]), .ready(ctrl_bus[5]), 
    .addr_(), .wdata(vga_cursor_wdata), .rdata(vga_cursor_rdata), 
	 .r_(vga_cursor_r), .w_(vga_cursor_w), .ready_(1'b1)
    );
wire [31:0]vga_text_addr, vga_text_wdata, vga_text_rdata;
wire vga_text_r;
wire [3:0]vga_text_w;
bus_interface VGA_TEXT(
    .enable(en_textRAM), 
    .addr(addr_bus), .data(data_bus), .r(ctrl_bus[0]), .w(ctrl_bus[4:1]), .ready(ctrl_bus[5]), 
    .addr_(vga_text_addr), .wdata(vga_text_wdata), .rdata(vga_text_rdata), 
	 .r_(vga_text_r), .w_(vga_text_w), .ready_(1'b1)
    );
wire [31:0]vga_graph_addr, vga_graph_wdata, vga_graph_rdata;
wire vga_graph_r;
wire [3:0]vga_graph_w;
bus_interface VGA_GRAPH(
    .enable(en_graphRAM), 
    .addr(addr_bus), .data(data_bus), .r(ctrl_bus[0]), .w(ctrl_bus[4:1]), .ready(ctrl_bus[5]), 
    .addr_(vga_graph_addr), .wdata(vga_graph_wdata), .rdata(vga_graph_rdata), 
	 .r_(vga_graph_r), .w_(vga_graph_w), .ready_(1'b1)
    );
wire SEG_r;
wire [3:0]SEG_w;
wire [31:0]SEG_wdata;
bus_interface SEG(
    .enable(en_SEG), 
    .addr(addr_bus), .data(data_bus), .r(ctrl_bus[0]), .w(ctrl_bus[4:1]), .ready(ctrl_bus[5]), 
    .addr_(), .wdata(SEG_wdata), .rdata(32'h0), 
	 .r_(SEG_r), .w_(SEG_w), .ready_(1'b1)
    );
wire keyboard_r;
wire [7:0]keyboard_data;
bus_interface keyboard(
    .enable(en_keyboard), 
    .addr(addr_bus), .data(data_bus), .r(ctrl_bus[0]), .w(ctrl_bus[4:1]), .ready(ctrl_bus[5]), 
    .addr_(), .wdata(), .rdata({24'b0, keyboard_data}),
	 .r_(keyboard_r), .w_(), .ready_(1'b1)
    );
bus_interface SWITCH(
    .enable(en_switch), 
    .addr(addr_bus), .data(data_bus), .r(ctrl_bus[0]), .w(ctrl_bus[4:1]), .ready(ctrl_bus[5]), 
    .addr_(), .wdata(), .rdata({16'b0, SW_OK[15:0]}), 
	 .r_(), .w_(), .ready_(1'b1)
    );
wire led_r;
wire [3:0]led_w;
wire [31:0]led_wdata, led_rdata;
bus_interface led(
    .enable(en_led), 
    .addr(addr_bus), .data(data_bus), .r(ctrl_bus[0]), .w(ctrl_bus[4:1]), .ready(ctrl_bus[5]), 
    .addr_(), .wdata(led_wdata), .rdata(led_rdata), 
	 .r_(led_r), .w_(led_w), .ready_(1'b1)
    );
wire dma_r;
wire [3:0]dma_w;
wire [31:0]dma_wdata, dma_rdata;
bus_interface dma(
    .enable(en_dma), 
    .addr(addr_bus), .data(data_bus), .r(ctrl_bus[0]), .w(ctrl_bus[4:1]), .ready(ctrl_bus[5]), 
    .addr_(), .wdata(dma_wdata), .rdata(dma_rdata), 
	 .r_(dma_r), .w_(dma_w), .ready_(1'b1)
    );
wire dmaRAM_r;
wire [3:0]dmaRAM_w;
wire [31:0]dmaRAM_wdata, dmaRAM_rdata;
wire [31:0]dmaRAM_addr;
bus_interface dmaRAM(
    .enable(en_dmaRAM), 
    .addr(addr_bus), .data(data_bus), .r(ctrl_bus[0]), .w(ctrl_bus[4:1]), .ready(ctrl_bus[5]), 
    .addr_(dmaRAM_addr), .wdata(dmaRAM_wdata), .rdata(dmaRAM_rdata), 
	 .r_(dmaRAM_r), .w_(dmaRAM_w), .ready_(1'b1)
    );
	 
wire [31:0]Disp_num;
wire [7:0]point_out;
wire [7:0]LE_out;
	 Display display(
    .clk(clk_100mhz), 
    .rst(rst), 
    .Start(Div[20]), 
    .Text(SW_OK[0]), 
    .flash(Div[25]), 
    .Hexs(Disp_num), 
    .point(point_out), 
    .LES(LE_out), 
    .segclk(seg_clk), 
    .segsout(seg_do), 
    .SEGEN(seg_pen), 
    .segclrn()
    );

wire [31:0]PC;
wire [31:0]inst;
wire [31:0]Data_in;
wire [31:0]cause_data;
wire [31:0]status_data;
wire [31:0]epc_data;
	Multi_8CH32  multi_8ch32(
		.clk(~Clk_CPU), 
		.Data0(SEG_wdata), 
		.data1(cause_data[31:0]), 
		.data2(inst[31:0]), 
		.data3(status_data[31:0]), 
		.data4(addr_bus[31:0]), 
		.data5(data_bus[31:0]), 
		.data6(epc_data[31:0]),
		.data7(PC[31:0]), 
		.EN(SEG_w), 
		.LES(64'b0), 
		.point_in({Div[31:0], Div[31:0]}), 
		.rst(rst), 
		.Test(SW_OK[7:5]), 
		.Disp_num(Disp_num), 
		.LE_out(LE_out), 
		.point_out(point_out)
		);

vga_controller Vga_controller(
    .clk(clk_100mhz), 
    .rst(rst), 
    .clk_vga(Div[1]), 
    .clk_cursor(Div[25]), 
    .we_text(vga_text_w), 
    .we_graph(vga_graph_w), 
    .we_cursor(vga_cursor_w), 
    .we_reg(vga_reg_w), 
	 .rd_text(vga_text_r), 
    .rd_graph(vga_graph_r), 
    .rd_cursor(vga_cursor_r), 
    .rd_reg(vga_reg_r), 
    .text_addr(vga_text_addr), 
    .text_wdata(vga_text_wdata), 
    .text_rdata(vga_text_rdata), 
    .graph_addr(vga_graph_addr), 
    .graph_wdata(vga_graph_wdata), 
    .graph_rdata(vga_graph_rdata), 
    .cursor_wdata(vga_cursor_wdata), 
    .cursor_rdata(vga_cursor_rdata), 
    .reg_wdata(vga_reg_wdata), 
    .reg_rdata(vga_reg_rdata), 
    .r(vga_red), 
    .g(vga_green), 
    .b(vga_blue), 
    .hsync(vga_h_sync), 
    .vsync(vga_v_sync), 
    .busy()
    );

wire keyboard_int;
keyboard_controller Keyboard_controller(
    .clk(clk_100mhz), 
    .clk_read(Clk_CPU),
    .rst(rst), 
    .ps2_clk(ps2_clk), 
    .ps2_data(ps2_dat), 
    .read(keyboard_r), 
    .ready(keyboard_int), 
    .full(), 
    .key_out(keyboard_data)
    );

led_controller Led_controller(
    .clk(clk_100mhz), 
    .rst(rst), 
    .we(led_w), 
    .wdata(led_wdata), 
    .rdata(led_rdata), 
    .led_clk(led_clk), 
    .led_do(led_do), 
    .led_pen(led_pen)
    );
	 
wire [31:0]CPU_wdata;
wire [31:0]CPU_mem_addr;
   PCPU_v PCPU(
		.clk(Clk_CPU), 
		`ifdef DEBUG
		.rst(RSTN),
		.int_(int_),
		`else
		.rst(rst),
		.int_({keyboard_int, 4'b0}),
		`endif
		.mem_we(ctrl_bus[4:1]), 
		.mem_rd(ctrl_bus[0]),
		.mem_addr(CPU_mem_addr), 
		.mem_data(CPU_wdata), 
		.inst_addr(PC), 
		.inst_data(inst), 
		.cause_data(cause_data),
		.status_data(status_data),
		.epc_data(epc_data),
		.mem_data_in(data_bus)
   );
assign addr_bus = {3'b0, CPU_mem_addr[28:0]};
assign data_bus = (|ctrl_bus[4:1]) ? CPU_wdata : 32'hz;
	/*
	Data_RAM Data_RAM_(
	  .clka(~Clk_CPU), 
	  .wea(SRAM_w), 
	  .addra(SRAM_addr[11:2]), 
	  .dina(SRAM_wdata), 
	  .douta(SRAM_rdata) 
	);
	*/
	wire [31:0]instBIOS;
	Inst_ROM BIOS(
	  .clka(~Clk_CPU), 
	  .addra(PC[11:2]), // addra,Ҫ�ƶ���λ
	  .douta(instBIOS) 
	);
	
	wire [31:0]instText;
	Text_Section TEXT(
  .clka(~Clk_CPU), 
  .wea(4'b0), 
  .addra(PC[12:2]), 
  .dina(32'b0), 
  .douta(instText), 
  .clkb(~Clk_CPU), 
  .web(TEXTS_bw), 
  .addrb(TEXTS_baddr), 
  .dinb(TEXTS_bwdata), 
  .doutb(TEXTS_brdata) 
  );
  assign inst = (PC[31:28] == 4'h1)? instBIOS : instText;

Data_Section DATA(
  .clka(~Clk_CPU), 
  .wea(DATAS_bw), 
  .addra(DATAS_baddr[31:2]), 
  .dina(DATAS_bwdata), 
  .douta(DATAS_brdata) 
);

/////////////////////////////////////////////////////
//DMA
wire [3:0]dma_mem_we;
wire [31:0]dma_mem_addr;
wire [31:0]dma_mem_rdata, dma_mem_wdata;
uart_controller UART_ctrl(
    .clk(clk_100mhz),
	 .clk_CPU(Clk_CPU),
    .rst(rst), 
    .we(dma_w),
    .rd(dma_r),
    .wdata(dma_wdata),
    .status(dma_rdata),  
    .mem_we(dma_mem_we), 
    .mem_addr(dma_mem_addr), 
    .mem_rdata(dma_mem_rdata), 
    .mem_wdata(dma_mem_wdata), 
    .rx_in(uart_rx), 
    .tx_out(uart_tx)
    );
	 
DMA_RAM DMA_RAM_(
  .clka(~Clk_CPU), // input clka
  .wea(dmaRAM_w), // input [3 : 0] wea
  .addra(dmaRAM_addr[8:2]), // input [6 : 0] addra
  .dina(dmaRAM_wdata), // input [31 : 0] dina
  .douta(dmaRAM_rdata), // output [31 : 0] douta
  .clkb(clk_100mhz), // input clkb
  .web(dma_mem_we), // input [3 : 0] web
  .addrb(dma_mem_addr[8:2]), // input [6 : 0] addrb
  .dinb(dma_mem_wdata), // input [31 : 0] dinb
  .doutb(dma_mem_rdata) // output [31 : 0] doutb
);

endmodule
