//`define DEBUG