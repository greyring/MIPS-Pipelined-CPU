`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    08:11:20 09/13/2017 
// Design Name: 
// Module Name:    mul32 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module mulu32(
	input [31:0]A,
	input [31:0]B,
	output [63:0]C
    );

wire c1_1_1, s1_1_1;
half_adder ha1_1_1 (
.a(A[0] & B[1]),.b(A[1] & B[0]),.p(s1_1_1),.g(c1_1_1)
);
wire c1_2_1, s1_2_1;
full_adder fa1_2_1 (
.a(A[0] & B[2]),.b(A[1] & B[1]),.c(A[2] & B[0]),.s(s1_2_1),.co(c1_2_1)
);
wire c1_3_1, s1_3_1;
full_adder fa1_3_1 (
.a(A[0] & B[3]),.b(A[1] & B[2]),.c(A[2] & B[1]),.s(s1_3_1),.co(c1_3_1)
);
wire c1_4_1, s1_4_1;
full_adder fa1_4_1 (
.a(A[0] & B[4]),.b(A[1] & B[3]),.c(A[2] & B[2]),.s(s1_4_1),.co(c1_4_1)
);
wire c1_4_2, s1_4_2;
half_adder ha1_4_2 (
.a(A[3] & B[1]),.b(A[4] & B[0]),.p(s1_4_2),.g(c1_4_2)
);
wire c1_5_1, s1_5_1;
full_adder fa1_5_1 (
.a(A[0] & B[5]),.b(A[1] & B[4]),.c(A[2] & B[3]),.s(s1_5_1),.co(c1_5_1)
);
wire c1_5_2, s1_5_2;
full_adder fa1_5_2 (
.a(A[3] & B[2]),.b(A[4] & B[1]),.c(A[5] & B[0]),.s(s1_5_2),.co(c1_5_2)
);
wire c1_6_1, s1_6_1;
full_adder fa1_6_1 (
.a(A[0] & B[6]),.b(A[1] & B[5]),.c(A[2] & B[4]),.s(s1_6_1),.co(c1_6_1)
);
wire c1_6_2, s1_6_2;
full_adder fa1_6_2 (
.a(A[3] & B[3]),.b(A[4] & B[2]),.c(A[5] & B[1]),.s(s1_6_2),.co(c1_6_2)
);
wire c1_7_1, s1_7_1;
full_adder fa1_7_1 (
.a(A[0] & B[7]),.b(A[1] & B[6]),.c(A[2] & B[5]),.s(s1_7_1),.co(c1_7_1)
);
wire c1_7_2, s1_7_2;
full_adder fa1_7_2 (
.a(A[3] & B[4]),.b(A[4] & B[3]),.c(A[5] & B[2]),.s(s1_7_2),.co(c1_7_2)
);
wire c1_7_3, s1_7_3;
half_adder ha1_7_3 (
.a(A[6] & B[1]),.b(A[7] & B[0]),.p(s1_7_3),.g(c1_7_3)
);
wire c1_8_1, s1_8_1;
full_adder fa1_8_1 (
.a(A[0] & B[8]),.b(A[1] & B[7]),.c(A[2] & B[6]),.s(s1_8_1),.co(c1_8_1)
);
wire c1_8_2, s1_8_2;
full_adder fa1_8_2 (
.a(A[3] & B[5]),.b(A[4] & B[4]),.c(A[5] & B[3]),.s(s1_8_2),.co(c1_8_2)
);
wire c1_8_3, s1_8_3;
full_adder fa1_8_3 (
.a(A[6] & B[2]),.b(A[7] & B[1]),.c(A[8] & B[0]),.s(s1_8_3),.co(c1_8_3)
);
wire c1_9_1, s1_9_1;
full_adder fa1_9_1 (
.a(A[0] & B[9]),.b(A[1] & B[8]),.c(A[2] & B[7]),.s(s1_9_1),.co(c1_9_1)
);
wire c1_9_2, s1_9_2;
full_adder fa1_9_2 (
.a(A[3] & B[6]),.b(A[4] & B[5]),.c(A[5] & B[4]),.s(s1_9_2),.co(c1_9_2)
);
wire c1_9_3, s1_9_3;
full_adder fa1_9_3 (
.a(A[6] & B[3]),.b(A[7] & B[2]),.c(A[8] & B[1]),.s(s1_9_3),.co(c1_9_3)
);
wire c1_10_1, s1_10_1;
full_adder fa1_10_1 (
.a(A[0] & B[10]),.b(A[1] & B[9]),.c(A[2] & B[8]),.s(s1_10_1),.co(c1_10_1)
);
wire c1_10_2, s1_10_2;
full_adder fa1_10_2 (
.a(A[3] & B[7]),.b(A[4] & B[6]),.c(A[5] & B[5]),.s(s1_10_2),.co(c1_10_2)
);
wire c1_10_3, s1_10_3;
full_adder fa1_10_3 (
.a(A[6] & B[4]),.b(A[7] & B[3]),.c(A[8] & B[2]),.s(s1_10_3),.co(c1_10_3)
);
wire c1_10_4, s1_10_4;
half_adder ha1_10_4 (
.a(A[9] & B[1]),.b(A[10] & B[0]),.p(s1_10_4),.g(c1_10_4)
);
wire c1_11_1, s1_11_1;
full_adder fa1_11_1 (
.a(A[0] & B[11]),.b(A[1] & B[10]),.c(A[2] & B[9]),.s(s1_11_1),.co(c1_11_1)
);
wire c1_11_2, s1_11_2;
full_adder fa1_11_2 (
.a(A[3] & B[8]),.b(A[4] & B[7]),.c(A[5] & B[6]),.s(s1_11_2),.co(c1_11_2)
);
wire c1_11_3, s1_11_3;
full_adder fa1_11_3 (
.a(A[6] & B[5]),.b(A[7] & B[4]),.c(A[8] & B[3]),.s(s1_11_3),.co(c1_11_3)
);
wire c1_11_4, s1_11_4;
full_adder fa1_11_4 (
.a(A[9] & B[2]),.b(A[10] & B[1]),.c(A[11] & B[0]),.s(s1_11_4),.co(c1_11_4)
);
wire c1_12_1, s1_12_1;
full_adder fa1_12_1 (
.a(A[0] & B[12]),.b(A[1] & B[11]),.c(A[2] & B[10]),.s(s1_12_1),.co(c1_12_1)
);
wire c1_12_2, s1_12_2;
full_adder fa1_12_2 (
.a(A[3] & B[9]),.b(A[4] & B[8]),.c(A[5] & B[7]),.s(s1_12_2),.co(c1_12_2)
);
wire c1_12_3, s1_12_3;
full_adder fa1_12_3 (
.a(A[6] & B[6]),.b(A[7] & B[5]),.c(A[8] & B[4]),.s(s1_12_3),.co(c1_12_3)
);
wire c1_12_4, s1_12_4;
full_adder fa1_12_4 (
.a(A[9] & B[3]),.b(A[10] & B[2]),.c(A[11] & B[1]),.s(s1_12_4),.co(c1_12_4)
);
wire c1_13_1, s1_13_1;
full_adder fa1_13_1 (
.a(A[0] & B[13]),.b(A[1] & B[12]),.c(A[2] & B[11]),.s(s1_13_1),.co(c1_13_1)
);
wire c1_13_2, s1_13_2;
full_adder fa1_13_2 (
.a(A[3] & B[10]),.b(A[4] & B[9]),.c(A[5] & B[8]),.s(s1_13_2),.co(c1_13_2)
);
wire c1_13_3, s1_13_3;
full_adder fa1_13_3 (
.a(A[6] & B[7]),.b(A[7] & B[6]),.c(A[8] & B[5]),.s(s1_13_3),.co(c1_13_3)
);
wire c1_13_4, s1_13_4;
full_adder fa1_13_4 (
.a(A[9] & B[4]),.b(A[10] & B[3]),.c(A[11] & B[2]),.s(s1_13_4),.co(c1_13_4)
);
wire c1_13_5, s1_13_5;
half_adder ha1_13_5 (
.a(A[12] & B[1]),.b(A[13] & B[0]),.p(s1_13_5),.g(c1_13_5)
);
wire c1_14_1, s1_14_1;
full_adder fa1_14_1 (
.a(A[0] & B[14]),.b(A[1] & B[13]),.c(A[2] & B[12]),.s(s1_14_1),.co(c1_14_1)
);
wire c1_14_2, s1_14_2;
full_adder fa1_14_2 (
.a(A[3] & B[11]),.b(A[4] & B[10]),.c(A[5] & B[9]),.s(s1_14_2),.co(c1_14_2)
);
wire c1_14_3, s1_14_3;
full_adder fa1_14_3 (
.a(A[6] & B[8]),.b(A[7] & B[7]),.c(A[8] & B[6]),.s(s1_14_3),.co(c1_14_3)
);
wire c1_14_4, s1_14_4;
full_adder fa1_14_4 (
.a(A[9] & B[5]),.b(A[10] & B[4]),.c(A[11] & B[3]),.s(s1_14_4),.co(c1_14_4)
);
wire c1_14_5, s1_14_5;
full_adder fa1_14_5 (
.a(A[12] & B[2]),.b(A[13] & B[1]),.c(A[14] & B[0]),.s(s1_14_5),.co(c1_14_5)
);
wire c1_15_1, s1_15_1;
full_adder fa1_15_1 (
.a(A[0] & B[15]),.b(A[1] & B[14]),.c(A[2] & B[13]),.s(s1_15_1),.co(c1_15_1)
);
wire c1_15_2, s1_15_2;
full_adder fa1_15_2 (
.a(A[3] & B[12]),.b(A[4] & B[11]),.c(A[5] & B[10]),.s(s1_15_2),.co(c1_15_2)
);
wire c1_15_3, s1_15_3;
full_adder fa1_15_3 (
.a(A[6] & B[9]),.b(A[7] & B[8]),.c(A[8] & B[7]),.s(s1_15_3),.co(c1_15_3)
);
wire c1_15_4, s1_15_4;
full_adder fa1_15_4 (
.a(A[9] & B[6]),.b(A[10] & B[5]),.c(A[11] & B[4]),.s(s1_15_4),.co(c1_15_4)
);
wire c1_15_5, s1_15_5;
full_adder fa1_15_5 (
.a(A[12] & B[3]),.b(A[13] & B[2]),.c(A[14] & B[1]),.s(s1_15_5),.co(c1_15_5)
);
wire c1_16_1, s1_16_1;
full_adder fa1_16_1 (
.a(A[0] & B[16]),.b(A[1] & B[15]),.c(A[2] & B[14]),.s(s1_16_1),.co(c1_16_1)
);
wire c1_16_2, s1_16_2;
full_adder fa1_16_2 (
.a(A[3] & B[13]),.b(A[4] & B[12]),.c(A[5] & B[11]),.s(s1_16_2),.co(c1_16_2)
);
wire c1_16_3, s1_16_3;
full_adder fa1_16_3 (
.a(A[6] & B[10]),.b(A[7] & B[9]),.c(A[8] & B[8]),.s(s1_16_3),.co(c1_16_3)
);
wire c1_16_4, s1_16_4;
full_adder fa1_16_4 (
.a(A[9] & B[7]),.b(A[10] & B[6]),.c(A[11] & B[5]),.s(s1_16_4),.co(c1_16_4)
);
wire c1_16_5, s1_16_5;
full_adder fa1_16_5 (
.a(A[12] & B[4]),.b(A[13] & B[3]),.c(A[14] & B[2]),.s(s1_16_5),.co(c1_16_5)
);
wire c1_16_6, s1_16_6;
half_adder ha1_16_6 (
.a(A[15] & B[1]),.b(A[16] & B[0]),.p(s1_16_6),.g(c1_16_6)
);
wire c1_17_1, s1_17_1;
full_adder fa1_17_1 (
.a(A[0] & B[17]),.b(A[1] & B[16]),.c(A[2] & B[15]),.s(s1_17_1),.co(c1_17_1)
);
wire c1_17_2, s1_17_2;
full_adder fa1_17_2 (
.a(A[3] & B[14]),.b(A[4] & B[13]),.c(A[5] & B[12]),.s(s1_17_2),.co(c1_17_2)
);
wire c1_17_3, s1_17_3;
full_adder fa1_17_3 (
.a(A[6] & B[11]),.b(A[7] & B[10]),.c(A[8] & B[9]),.s(s1_17_3),.co(c1_17_3)
);
wire c1_17_4, s1_17_4;
full_adder fa1_17_4 (
.a(A[9] & B[8]),.b(A[10] & B[7]),.c(A[11] & B[6]),.s(s1_17_4),.co(c1_17_4)
);
wire c1_17_5, s1_17_5;
full_adder fa1_17_5 (
.a(A[12] & B[5]),.b(A[13] & B[4]),.c(A[14] & B[3]),.s(s1_17_5),.co(c1_17_5)
);
wire c1_17_6, s1_17_6;
full_adder fa1_17_6 (
.a(A[15] & B[2]),.b(A[16] & B[1]),.c(A[17] & B[0]),.s(s1_17_6),.co(c1_17_6)
);
wire c1_18_1, s1_18_1;
full_adder fa1_18_1 (
.a(A[0] & B[18]),.b(A[1] & B[17]),.c(A[2] & B[16]),.s(s1_18_1),.co(c1_18_1)
);
wire c1_18_2, s1_18_2;
full_adder fa1_18_2 (
.a(A[3] & B[15]),.b(A[4] & B[14]),.c(A[5] & B[13]),.s(s1_18_2),.co(c1_18_2)
);
wire c1_18_3, s1_18_3;
full_adder fa1_18_3 (
.a(A[6] & B[12]),.b(A[7] & B[11]),.c(A[8] & B[10]),.s(s1_18_3),.co(c1_18_3)
);
wire c1_18_4, s1_18_4;
full_adder fa1_18_4 (
.a(A[9] & B[9]),.b(A[10] & B[8]),.c(A[11] & B[7]),.s(s1_18_4),.co(c1_18_4)
);
wire c1_18_5, s1_18_5;
full_adder fa1_18_5 (
.a(A[12] & B[6]),.b(A[13] & B[5]),.c(A[14] & B[4]),.s(s1_18_5),.co(c1_18_5)
);
wire c1_18_6, s1_18_6;
full_adder fa1_18_6 (
.a(A[15] & B[3]),.b(A[16] & B[2]),.c(A[17] & B[1]),.s(s1_18_6),.co(c1_18_6)
);
wire c1_19_1, s1_19_1;
full_adder fa1_19_1 (
.a(A[0] & B[19]),.b(A[1] & B[18]),.c(A[2] & B[17]),.s(s1_19_1),.co(c1_19_1)
);
wire c1_19_2, s1_19_2;
full_adder fa1_19_2 (
.a(A[3] & B[16]),.b(A[4] & B[15]),.c(A[5] & B[14]),.s(s1_19_2),.co(c1_19_2)
);
wire c1_19_3, s1_19_3;
full_adder fa1_19_3 (
.a(A[6] & B[13]),.b(A[7] & B[12]),.c(A[8] & B[11]),.s(s1_19_3),.co(c1_19_3)
);
wire c1_19_4, s1_19_4;
full_adder fa1_19_4 (
.a(A[9] & B[10]),.b(A[10] & B[9]),.c(A[11] & B[8]),.s(s1_19_4),.co(c1_19_4)
);
wire c1_19_5, s1_19_5;
full_adder fa1_19_5 (
.a(A[12] & B[7]),.b(A[13] & B[6]),.c(A[14] & B[5]),.s(s1_19_5),.co(c1_19_5)
);
wire c1_19_6, s1_19_6;
full_adder fa1_19_6 (
.a(A[15] & B[4]),.b(A[16] & B[3]),.c(A[17] & B[2]),.s(s1_19_6),.co(c1_19_6)
);
wire c1_19_7, s1_19_7;
half_adder ha1_19_7 (
.a(A[18] & B[1]),.b(A[19] & B[0]),.p(s1_19_7),.g(c1_19_7)
);
wire c1_20_1, s1_20_1;
full_adder fa1_20_1 (
.a(A[0] & B[20]),.b(A[1] & B[19]),.c(A[2] & B[18]),.s(s1_20_1),.co(c1_20_1)
);
wire c1_20_2, s1_20_2;
full_adder fa1_20_2 (
.a(A[3] & B[17]),.b(A[4] & B[16]),.c(A[5] & B[15]),.s(s1_20_2),.co(c1_20_2)
);
wire c1_20_3, s1_20_3;
full_adder fa1_20_3 (
.a(A[6] & B[14]),.b(A[7] & B[13]),.c(A[8] & B[12]),.s(s1_20_3),.co(c1_20_3)
);
wire c1_20_4, s1_20_4;
full_adder fa1_20_4 (
.a(A[9] & B[11]),.b(A[10] & B[10]),.c(A[11] & B[9]),.s(s1_20_4),.co(c1_20_4)
);
wire c1_20_5, s1_20_5;
full_adder fa1_20_5 (
.a(A[12] & B[8]),.b(A[13] & B[7]),.c(A[14] & B[6]),.s(s1_20_5),.co(c1_20_5)
);
wire c1_20_6, s1_20_6;
full_adder fa1_20_6 (
.a(A[15] & B[5]),.b(A[16] & B[4]),.c(A[17] & B[3]),.s(s1_20_6),.co(c1_20_6)
);
wire c1_20_7, s1_20_7;
full_adder fa1_20_7 (
.a(A[18] & B[2]),.b(A[19] & B[1]),.c(A[20] & B[0]),.s(s1_20_7),.co(c1_20_7)
);
wire c1_21_1, s1_21_1;
full_adder fa1_21_1 (
.a(A[0] & B[21]),.b(A[1] & B[20]),.c(A[2] & B[19]),.s(s1_21_1),.co(c1_21_1)
);
wire c1_21_2, s1_21_2;
full_adder fa1_21_2 (
.a(A[3] & B[18]),.b(A[4] & B[17]),.c(A[5] & B[16]),.s(s1_21_2),.co(c1_21_2)
);
wire c1_21_3, s1_21_3;
full_adder fa1_21_3 (
.a(A[6] & B[15]),.b(A[7] & B[14]),.c(A[8] & B[13]),.s(s1_21_3),.co(c1_21_3)
);
wire c1_21_4, s1_21_4;
full_adder fa1_21_4 (
.a(A[9] & B[12]),.b(A[10] & B[11]),.c(A[11] & B[10]),.s(s1_21_4),.co(c1_21_4)
);
wire c1_21_5, s1_21_5;
full_adder fa1_21_5 (
.a(A[12] & B[9]),.b(A[13] & B[8]),.c(A[14] & B[7]),.s(s1_21_5),.co(c1_21_5)
);
wire c1_21_6, s1_21_6;
full_adder fa1_21_6 (
.a(A[15] & B[6]),.b(A[16] & B[5]),.c(A[17] & B[4]),.s(s1_21_6),.co(c1_21_6)
);
wire c1_21_7, s1_21_7;
full_adder fa1_21_7 (
.a(A[18] & B[3]),.b(A[19] & B[2]),.c(A[20] & B[1]),.s(s1_21_7),.co(c1_21_7)
);
wire c1_22_1, s1_22_1;
full_adder fa1_22_1 (
.a(A[0] & B[22]),.b(A[1] & B[21]),.c(A[2] & B[20]),.s(s1_22_1),.co(c1_22_1)
);
wire c1_22_2, s1_22_2;
full_adder fa1_22_2 (
.a(A[3] & B[19]),.b(A[4] & B[18]),.c(A[5] & B[17]),.s(s1_22_2),.co(c1_22_2)
);
wire c1_22_3, s1_22_3;
full_adder fa1_22_3 (
.a(A[6] & B[16]),.b(A[7] & B[15]),.c(A[8] & B[14]),.s(s1_22_3),.co(c1_22_3)
);
wire c1_22_4, s1_22_4;
full_adder fa1_22_4 (
.a(A[9] & B[13]),.b(A[10] & B[12]),.c(A[11] & B[11]),.s(s1_22_4),.co(c1_22_4)
);
wire c1_22_5, s1_22_5;
full_adder fa1_22_5 (
.a(A[12] & B[10]),.b(A[13] & B[9]),.c(A[14] & B[8]),.s(s1_22_5),.co(c1_22_5)
);
wire c1_22_6, s1_22_6;
full_adder fa1_22_6 (
.a(A[15] & B[7]),.b(A[16] & B[6]),.c(A[17] & B[5]),.s(s1_22_6),.co(c1_22_6)
);
wire c1_22_7, s1_22_7;
full_adder fa1_22_7 (
.a(A[18] & B[4]),.b(A[19] & B[3]),.c(A[20] & B[2]),.s(s1_22_7),.co(c1_22_7)
);
wire c1_22_8, s1_22_8;
half_adder ha1_22_8 (
.a(A[21] & B[1]),.b(A[22] & B[0]),.p(s1_22_8),.g(c1_22_8)
);
wire c1_23_1, s1_23_1;
full_adder fa1_23_1 (
.a(A[0] & B[23]),.b(A[1] & B[22]),.c(A[2] & B[21]),.s(s1_23_1),.co(c1_23_1)
);
wire c1_23_2, s1_23_2;
full_adder fa1_23_2 (
.a(A[3] & B[20]),.b(A[4] & B[19]),.c(A[5] & B[18]),.s(s1_23_2),.co(c1_23_2)
);
wire c1_23_3, s1_23_3;
full_adder fa1_23_3 (
.a(A[6] & B[17]),.b(A[7] & B[16]),.c(A[8] & B[15]),.s(s1_23_3),.co(c1_23_3)
);
wire c1_23_4, s1_23_4;
full_adder fa1_23_4 (
.a(A[9] & B[14]),.b(A[10] & B[13]),.c(A[11] & B[12]),.s(s1_23_4),.co(c1_23_4)
);
wire c1_23_5, s1_23_5;
full_adder fa1_23_5 (
.a(A[12] & B[11]),.b(A[13] & B[10]),.c(A[14] & B[9]),.s(s1_23_5),.co(c1_23_5)
);
wire c1_23_6, s1_23_6;
full_adder fa1_23_6 (
.a(A[15] & B[8]),.b(A[16] & B[7]),.c(A[17] & B[6]),.s(s1_23_6),.co(c1_23_6)
);
wire c1_23_7, s1_23_7;
full_adder fa1_23_7 (
.a(A[18] & B[5]),.b(A[19] & B[4]),.c(A[20] & B[3]),.s(s1_23_7),.co(c1_23_7)
);
wire c1_23_8, s1_23_8;
full_adder fa1_23_8 (
.a(A[21] & B[2]),.b(A[22] & B[1]),.c(A[23] & B[0]),.s(s1_23_8),.co(c1_23_8)
);
wire c1_24_1, s1_24_1;
full_adder fa1_24_1 (
.a(A[0] & B[24]),.b(A[1] & B[23]),.c(A[2] & B[22]),.s(s1_24_1),.co(c1_24_1)
);
wire c1_24_2, s1_24_2;
full_adder fa1_24_2 (
.a(A[3] & B[21]),.b(A[4] & B[20]),.c(A[5] & B[19]),.s(s1_24_2),.co(c1_24_2)
);
wire c1_24_3, s1_24_3;
full_adder fa1_24_3 (
.a(A[6] & B[18]),.b(A[7] & B[17]),.c(A[8] & B[16]),.s(s1_24_3),.co(c1_24_3)
);
wire c1_24_4, s1_24_4;
full_adder fa1_24_4 (
.a(A[9] & B[15]),.b(A[10] & B[14]),.c(A[11] & B[13]),.s(s1_24_4),.co(c1_24_4)
);
wire c1_24_5, s1_24_5;
full_adder fa1_24_5 (
.a(A[12] & B[12]),.b(A[13] & B[11]),.c(A[14] & B[10]),.s(s1_24_5),.co(c1_24_5)
);
wire c1_24_6, s1_24_6;
full_adder fa1_24_6 (
.a(A[15] & B[9]),.b(A[16] & B[8]),.c(A[17] & B[7]),.s(s1_24_6),.co(c1_24_6)
);
wire c1_24_7, s1_24_7;
full_adder fa1_24_7 (
.a(A[18] & B[6]),.b(A[19] & B[5]),.c(A[20] & B[4]),.s(s1_24_7),.co(c1_24_7)
);
wire c1_24_8, s1_24_8;
full_adder fa1_24_8 (
.a(A[21] & B[3]),.b(A[22] & B[2]),.c(A[23] & B[1]),.s(s1_24_8),.co(c1_24_8)
);
wire c1_25_1, s1_25_1;
full_adder fa1_25_1 (
.a(A[0] & B[25]),.b(A[1] & B[24]),.c(A[2] & B[23]),.s(s1_25_1),.co(c1_25_1)
);
wire c1_25_2, s1_25_2;
full_adder fa1_25_2 (
.a(A[3] & B[22]),.b(A[4] & B[21]),.c(A[5] & B[20]),.s(s1_25_2),.co(c1_25_2)
);
wire c1_25_3, s1_25_3;
full_adder fa1_25_3 (
.a(A[6] & B[19]),.b(A[7] & B[18]),.c(A[8] & B[17]),.s(s1_25_3),.co(c1_25_3)
);
wire c1_25_4, s1_25_4;
full_adder fa1_25_4 (
.a(A[9] & B[16]),.b(A[10] & B[15]),.c(A[11] & B[14]),.s(s1_25_4),.co(c1_25_4)
);
wire c1_25_5, s1_25_5;
full_adder fa1_25_5 (
.a(A[12] & B[13]),.b(A[13] & B[12]),.c(A[14] & B[11]),.s(s1_25_5),.co(c1_25_5)
);
wire c1_25_6, s1_25_6;
full_adder fa1_25_6 (
.a(A[15] & B[10]),.b(A[16] & B[9]),.c(A[17] & B[8]),.s(s1_25_6),.co(c1_25_6)
);
wire c1_25_7, s1_25_7;
full_adder fa1_25_7 (
.a(A[18] & B[7]),.b(A[19] & B[6]),.c(A[20] & B[5]),.s(s1_25_7),.co(c1_25_7)
);
wire c1_25_8, s1_25_8;
full_adder fa1_25_8 (
.a(A[21] & B[4]),.b(A[22] & B[3]),.c(A[23] & B[2]),.s(s1_25_8),.co(c1_25_8)
);
wire c1_25_9, s1_25_9;
half_adder ha1_25_9 (
.a(A[24] & B[1]),.b(A[25] & B[0]),.p(s1_25_9),.g(c1_25_9)
);
wire c1_26_1, s1_26_1;
full_adder fa1_26_1 (
.a(A[0] & B[26]),.b(A[1] & B[25]),.c(A[2] & B[24]),.s(s1_26_1),.co(c1_26_1)
);
wire c1_26_2, s1_26_2;
full_adder fa1_26_2 (
.a(A[3] & B[23]),.b(A[4] & B[22]),.c(A[5] & B[21]),.s(s1_26_2),.co(c1_26_2)
);
wire c1_26_3, s1_26_3;
full_adder fa1_26_3 (
.a(A[6] & B[20]),.b(A[7] & B[19]),.c(A[8] & B[18]),.s(s1_26_3),.co(c1_26_3)
);
wire c1_26_4, s1_26_4;
full_adder fa1_26_4 (
.a(A[9] & B[17]),.b(A[10] & B[16]),.c(A[11] & B[15]),.s(s1_26_4),.co(c1_26_4)
);
wire c1_26_5, s1_26_5;
full_adder fa1_26_5 (
.a(A[12] & B[14]),.b(A[13] & B[13]),.c(A[14] & B[12]),.s(s1_26_5),.co(c1_26_5)
);
wire c1_26_6, s1_26_6;
full_adder fa1_26_6 (
.a(A[15] & B[11]),.b(A[16] & B[10]),.c(A[17] & B[9]),.s(s1_26_6),.co(c1_26_6)
);
wire c1_26_7, s1_26_7;
full_adder fa1_26_7 (
.a(A[18] & B[8]),.b(A[19] & B[7]),.c(A[20] & B[6]),.s(s1_26_7),.co(c1_26_7)
);
wire c1_26_8, s1_26_8;
full_adder fa1_26_8 (
.a(A[21] & B[5]),.b(A[22] & B[4]),.c(A[23] & B[3]),.s(s1_26_8),.co(c1_26_8)
);
wire c1_26_9, s1_26_9;
full_adder fa1_26_9 (
.a(A[24] & B[2]),.b(A[25] & B[1]),.c(A[26] & B[0]),.s(s1_26_9),.co(c1_26_9)
);
wire c1_27_1, s1_27_1;
full_adder fa1_27_1 (
.a(A[0] & B[27]),.b(A[1] & B[26]),.c(A[2] & B[25]),.s(s1_27_1),.co(c1_27_1)
);
wire c1_27_2, s1_27_2;
full_adder fa1_27_2 (
.a(A[3] & B[24]),.b(A[4] & B[23]),.c(A[5] & B[22]),.s(s1_27_2),.co(c1_27_2)
);
wire c1_27_3, s1_27_3;
full_adder fa1_27_3 (
.a(A[6] & B[21]),.b(A[7] & B[20]),.c(A[8] & B[19]),.s(s1_27_3),.co(c1_27_3)
);
wire c1_27_4, s1_27_4;
full_adder fa1_27_4 (
.a(A[9] & B[18]),.b(A[10] & B[17]),.c(A[11] & B[16]),.s(s1_27_4),.co(c1_27_4)
);
wire c1_27_5, s1_27_5;
full_adder fa1_27_5 (
.a(A[12] & B[15]),.b(A[13] & B[14]),.c(A[14] & B[13]),.s(s1_27_5),.co(c1_27_5)
);
wire c1_27_6, s1_27_6;
full_adder fa1_27_6 (
.a(A[15] & B[12]),.b(A[16] & B[11]),.c(A[17] & B[10]),.s(s1_27_6),.co(c1_27_6)
);
wire c1_27_7, s1_27_7;
full_adder fa1_27_7 (
.a(A[18] & B[9]),.b(A[19] & B[8]),.c(A[20] & B[7]),.s(s1_27_7),.co(c1_27_7)
);
wire c1_27_8, s1_27_8;
full_adder fa1_27_8 (
.a(A[21] & B[6]),.b(A[22] & B[5]),.c(A[23] & B[4]),.s(s1_27_8),.co(c1_27_8)
);
wire c1_27_9, s1_27_9;
full_adder fa1_27_9 (
.a(A[24] & B[3]),.b(A[25] & B[2]),.c(A[26] & B[1]),.s(s1_27_9),.co(c1_27_9)
);
wire c1_28_1, s1_28_1;
full_adder fa1_28_1 (
.a(A[0] & B[28]),.b(A[1] & B[27]),.c(A[2] & B[26]),.s(s1_28_1),.co(c1_28_1)
);
wire c1_28_2, s1_28_2;
full_adder fa1_28_2 (
.a(A[3] & B[25]),.b(A[4] & B[24]),.c(A[5] & B[23]),.s(s1_28_2),.co(c1_28_2)
);
wire c1_28_3, s1_28_3;
full_adder fa1_28_3 (
.a(A[6] & B[22]),.b(A[7] & B[21]),.c(A[8] & B[20]),.s(s1_28_3),.co(c1_28_3)
);
wire c1_28_4, s1_28_4;
full_adder fa1_28_4 (
.a(A[9] & B[19]),.b(A[10] & B[18]),.c(A[11] & B[17]),.s(s1_28_4),.co(c1_28_4)
);
wire c1_28_5, s1_28_5;
full_adder fa1_28_5 (
.a(A[12] & B[16]),.b(A[13] & B[15]),.c(A[14] & B[14]),.s(s1_28_5),.co(c1_28_5)
);
wire c1_28_6, s1_28_6;
full_adder fa1_28_6 (
.a(A[15] & B[13]),.b(A[16] & B[12]),.c(A[17] & B[11]),.s(s1_28_6),.co(c1_28_6)
);
wire c1_28_7, s1_28_7;
full_adder fa1_28_7 (
.a(A[18] & B[10]),.b(A[19] & B[9]),.c(A[20] & B[8]),.s(s1_28_7),.co(c1_28_7)
);
wire c1_28_8, s1_28_8;
full_adder fa1_28_8 (
.a(A[21] & B[7]),.b(A[22] & B[6]),.c(A[23] & B[5]),.s(s1_28_8),.co(c1_28_8)
);
wire c1_28_9, s1_28_9;
full_adder fa1_28_9 (
.a(A[24] & B[4]),.b(A[25] & B[3]),.c(A[26] & B[2]),.s(s1_28_9),.co(c1_28_9)
);
wire c1_28_10, s1_28_10;
half_adder ha1_28_10 (
.a(A[27] & B[1]),.b(A[28] & B[0]),.p(s1_28_10),.g(c1_28_10)
);
wire c1_29_1, s1_29_1;
full_adder fa1_29_1 (
.a(A[0] & B[29]),.b(A[1] & B[28]),.c(A[2] & B[27]),.s(s1_29_1),.co(c1_29_1)
);
wire c1_29_2, s1_29_2;
full_adder fa1_29_2 (
.a(A[3] & B[26]),.b(A[4] & B[25]),.c(A[5] & B[24]),.s(s1_29_2),.co(c1_29_2)
);
wire c1_29_3, s1_29_3;
full_adder fa1_29_3 (
.a(A[6] & B[23]),.b(A[7] & B[22]),.c(A[8] & B[21]),.s(s1_29_3),.co(c1_29_3)
);
wire c1_29_4, s1_29_4;
full_adder fa1_29_4 (
.a(A[9] & B[20]),.b(A[10] & B[19]),.c(A[11] & B[18]),.s(s1_29_4),.co(c1_29_4)
);
wire c1_29_5, s1_29_5;
full_adder fa1_29_5 (
.a(A[12] & B[17]),.b(A[13] & B[16]),.c(A[14] & B[15]),.s(s1_29_5),.co(c1_29_5)
);
wire c1_29_6, s1_29_6;
full_adder fa1_29_6 (
.a(A[15] & B[14]),.b(A[16] & B[13]),.c(A[17] & B[12]),.s(s1_29_6),.co(c1_29_6)
);
wire c1_29_7, s1_29_7;
full_adder fa1_29_7 (
.a(A[18] & B[11]),.b(A[19] & B[10]),.c(A[20] & B[9]),.s(s1_29_7),.co(c1_29_7)
);
wire c1_29_8, s1_29_8;
full_adder fa1_29_8 (
.a(A[21] & B[8]),.b(A[22] & B[7]),.c(A[23] & B[6]),.s(s1_29_8),.co(c1_29_8)
);
wire c1_29_9, s1_29_9;
full_adder fa1_29_9 (
.a(A[24] & B[5]),.b(A[25] & B[4]),.c(A[26] & B[3]),.s(s1_29_9),.co(c1_29_9)
);
wire c1_29_10, s1_29_10;
full_adder fa1_29_10 (
.a(A[27] & B[2]),.b(A[28] & B[1]),.c(A[29] & B[0]),.s(s1_29_10),.co(c1_29_10)
);
wire c1_30_1, s1_30_1;
full_adder fa1_30_1 (
.a(A[0] & B[30]),.b(A[1] & B[29]),.c(A[2] & B[28]),.s(s1_30_1),.co(c1_30_1)
);
wire c1_30_2, s1_30_2;
full_adder fa1_30_2 (
.a(A[3] & B[27]),.b(A[4] & B[26]),.c(A[5] & B[25]),.s(s1_30_2),.co(c1_30_2)
);
wire c1_30_3, s1_30_3;
full_adder fa1_30_3 (
.a(A[6] & B[24]),.b(A[7] & B[23]),.c(A[8] & B[22]),.s(s1_30_3),.co(c1_30_3)
);
wire c1_30_4, s1_30_4;
full_adder fa1_30_4 (
.a(A[9] & B[21]),.b(A[10] & B[20]),.c(A[11] & B[19]),.s(s1_30_4),.co(c1_30_4)
);
wire c1_30_5, s1_30_5;
full_adder fa1_30_5 (
.a(A[12] & B[18]),.b(A[13] & B[17]),.c(A[14] & B[16]),.s(s1_30_5),.co(c1_30_5)
);
wire c1_30_6, s1_30_6;
full_adder fa1_30_6 (
.a(A[15] & B[15]),.b(A[16] & B[14]),.c(A[17] & B[13]),.s(s1_30_6),.co(c1_30_6)
);
wire c1_30_7, s1_30_7;
full_adder fa1_30_7 (
.a(A[18] & B[12]),.b(A[19] & B[11]),.c(A[20] & B[10]),.s(s1_30_7),.co(c1_30_7)
);
wire c1_30_8, s1_30_8;
full_adder fa1_30_8 (
.a(A[21] & B[9]),.b(A[22] & B[8]),.c(A[23] & B[7]),.s(s1_30_8),.co(c1_30_8)
);
wire c1_30_9, s1_30_9;
full_adder fa1_30_9 (
.a(A[24] & B[6]),.b(A[25] & B[5]),.c(A[26] & B[4]),.s(s1_30_9),.co(c1_30_9)
);
wire c1_30_10, s1_30_10;
full_adder fa1_30_10 (
.a(A[27] & B[3]),.b(A[28] & B[2]),.c(A[29] & B[1]),.s(s1_30_10),.co(c1_30_10)
);
wire c1_31_1, s1_31_1;
full_adder fa1_31_1 (
.a(A[0] & B[31]),.b(A[1] & B[30]),.c(A[2] & B[29]),.s(s1_31_1),.co(c1_31_1)
);
wire c1_31_2, s1_31_2;
full_adder fa1_31_2 (
.a(A[3] & B[28]),.b(A[4] & B[27]),.c(A[5] & B[26]),.s(s1_31_2),.co(c1_31_2)
);
wire c1_31_3, s1_31_3;
full_adder fa1_31_3 (
.a(A[6] & B[25]),.b(A[7] & B[24]),.c(A[8] & B[23]),.s(s1_31_3),.co(c1_31_3)
);
wire c1_31_4, s1_31_4;
full_adder fa1_31_4 (
.a(A[9] & B[22]),.b(A[10] & B[21]),.c(A[11] & B[20]),.s(s1_31_4),.co(c1_31_4)
);
wire c1_31_5, s1_31_5;
full_adder fa1_31_5 (
.a(A[12] & B[19]),.b(A[13] & B[18]),.c(A[14] & B[17]),.s(s1_31_5),.co(c1_31_5)
);
wire c1_31_6, s1_31_6;
full_adder fa1_31_6 (
.a(A[15] & B[16]),.b(A[16] & B[15]),.c(A[17] & B[14]),.s(s1_31_6),.co(c1_31_6)
);
wire c1_31_7, s1_31_7;
full_adder fa1_31_7 (
.a(A[18] & B[13]),.b(A[19] & B[12]),.c(A[20] & B[11]),.s(s1_31_7),.co(c1_31_7)
);
wire c1_31_8, s1_31_8;
full_adder fa1_31_8 (
.a(A[21] & B[10]),.b(A[22] & B[9]),.c(A[23] & B[8]),.s(s1_31_8),.co(c1_31_8)
);
wire c1_31_9, s1_31_9;
full_adder fa1_31_9 (
.a(A[24] & B[7]),.b(A[25] & B[6]),.c(A[26] & B[5]),.s(s1_31_9),.co(c1_31_9)
);
wire c1_31_10, s1_31_10;
full_adder fa1_31_10 (
.a(A[27] & B[4]),.b(A[28] & B[3]),.c(A[29] & B[2]),.s(s1_31_10),.co(c1_31_10)
);
wire c1_31_11, s1_31_11;
half_adder ha1_31_11 (
.a(A[30] & B[1]),.b(A[31] & B[0]),.p(s1_31_11),.g(c1_31_11)
);
wire c1_32_1, s1_32_1;
full_adder fa1_32_1 (
.a(A[1] & B[31]),.b(A[2] & B[30]),.c(A[3] & B[29]),.s(s1_32_1),.co(c1_32_1)
);
wire c1_32_2, s1_32_2;
full_adder fa1_32_2 (
.a(A[4] & B[28]),.b(A[5] & B[27]),.c(A[6] & B[26]),.s(s1_32_2),.co(c1_32_2)
);
wire c1_32_3, s1_32_3;
full_adder fa1_32_3 (
.a(A[7] & B[25]),.b(A[8] & B[24]),.c(A[9] & B[23]),.s(s1_32_3),.co(c1_32_3)
);
wire c1_32_4, s1_32_4;
full_adder fa1_32_4 (
.a(A[10] & B[22]),.b(A[11] & B[21]),.c(A[12] & B[20]),.s(s1_32_4),.co(c1_32_4)
);
wire c1_32_5, s1_32_5;
full_adder fa1_32_5 (
.a(A[13] & B[19]),.b(A[14] & B[18]),.c(A[15] & B[17]),.s(s1_32_5),.co(c1_32_5)
);
wire c1_32_6, s1_32_6;
full_adder fa1_32_6 (
.a(A[16] & B[16]),.b(A[17] & B[15]),.c(A[18] & B[14]),.s(s1_32_6),.co(c1_32_6)
);
wire c1_32_7, s1_32_7;
full_adder fa1_32_7 (
.a(A[19] & B[13]),.b(A[20] & B[12]),.c(A[21] & B[11]),.s(s1_32_7),.co(c1_32_7)
);
wire c1_32_8, s1_32_8;
full_adder fa1_32_8 (
.a(A[22] & B[10]),.b(A[23] & B[9]),.c(A[24] & B[8]),.s(s1_32_8),.co(c1_32_8)
);
wire c1_32_9, s1_32_9;
full_adder fa1_32_9 (
.a(A[25] & B[7]),.b(A[26] & B[6]),.c(A[27] & B[5]),.s(s1_32_9),.co(c1_32_9)
);
wire c1_32_10, s1_32_10;
full_adder fa1_32_10 (
.a(A[28] & B[4]),.b(A[29] & B[3]),.c(A[30] & B[2]),.s(s1_32_10),.co(c1_32_10)
);
wire c1_33_1, s1_33_1;
full_adder fa1_33_1 (
.a(A[2] & B[31]),.b(A[3] & B[30]),.c(A[4] & B[29]),.s(s1_33_1),.co(c1_33_1)
);
wire c1_33_2, s1_33_2;
full_adder fa1_33_2 (
.a(A[5] & B[28]),.b(A[6] & B[27]),.c(A[7] & B[26]),.s(s1_33_2),.co(c1_33_2)
);
wire c1_33_3, s1_33_3;
full_adder fa1_33_3 (
.a(A[8] & B[25]),.b(A[9] & B[24]),.c(A[10] & B[23]),.s(s1_33_3),.co(c1_33_3)
);
wire c1_33_4, s1_33_4;
full_adder fa1_33_4 (
.a(A[11] & B[22]),.b(A[12] & B[21]),.c(A[13] & B[20]),.s(s1_33_4),.co(c1_33_4)
);
wire c1_33_5, s1_33_5;
full_adder fa1_33_5 (
.a(A[14] & B[19]),.b(A[15] & B[18]),.c(A[16] & B[17]),.s(s1_33_5),.co(c1_33_5)
);
wire c1_33_6, s1_33_6;
full_adder fa1_33_6 (
.a(A[17] & B[16]),.b(A[18] & B[15]),.c(A[19] & B[14]),.s(s1_33_6),.co(c1_33_6)
);
wire c1_33_7, s1_33_7;
full_adder fa1_33_7 (
.a(A[20] & B[13]),.b(A[21] & B[12]),.c(A[22] & B[11]),.s(s1_33_7),.co(c1_33_7)
);
wire c1_33_8, s1_33_8;
full_adder fa1_33_8 (
.a(A[23] & B[10]),.b(A[24] & B[9]),.c(A[25] & B[8]),.s(s1_33_8),.co(c1_33_8)
);
wire c1_33_9, s1_33_9;
full_adder fa1_33_9 (
.a(A[26] & B[7]),.b(A[27] & B[6]),.c(A[28] & B[5]),.s(s1_33_9),.co(c1_33_9)
);
wire c1_33_10, s1_33_10;
full_adder fa1_33_10 (
.a(A[29] & B[4]),.b(A[30] & B[3]),.c(A[31] & B[2]),.s(s1_33_10),.co(c1_33_10)
);
wire c1_34_1, s1_34_1;
full_adder fa1_34_1 (
.a(A[3] & B[31]),.b(A[4] & B[30]),.c(A[5] & B[29]),.s(s1_34_1),.co(c1_34_1)
);
wire c1_34_2, s1_34_2;
full_adder fa1_34_2 (
.a(A[6] & B[28]),.b(A[7] & B[27]),.c(A[8] & B[26]),.s(s1_34_2),.co(c1_34_2)
);
wire c1_34_3, s1_34_3;
full_adder fa1_34_3 (
.a(A[9] & B[25]),.b(A[10] & B[24]),.c(A[11] & B[23]),.s(s1_34_3),.co(c1_34_3)
);
wire c1_34_4, s1_34_4;
full_adder fa1_34_4 (
.a(A[12] & B[22]),.b(A[13] & B[21]),.c(A[14] & B[20]),.s(s1_34_4),.co(c1_34_4)
);
wire c1_34_5, s1_34_5;
full_adder fa1_34_5 (
.a(A[15] & B[19]),.b(A[16] & B[18]),.c(A[17] & B[17]),.s(s1_34_5),.co(c1_34_5)
);
wire c1_34_6, s1_34_6;
full_adder fa1_34_6 (
.a(A[18] & B[16]),.b(A[19] & B[15]),.c(A[20] & B[14]),.s(s1_34_6),.co(c1_34_6)
);
wire c1_34_7, s1_34_7;
full_adder fa1_34_7 (
.a(A[21] & B[13]),.b(A[22] & B[12]),.c(A[23] & B[11]),.s(s1_34_7),.co(c1_34_7)
);
wire c1_34_8, s1_34_8;
full_adder fa1_34_8 (
.a(A[24] & B[10]),.b(A[25] & B[9]),.c(A[26] & B[8]),.s(s1_34_8),.co(c1_34_8)
);
wire c1_34_9, s1_34_9;
full_adder fa1_34_9 (
.a(A[27] & B[7]),.b(A[28] & B[6]),.c(A[29] & B[5]),.s(s1_34_9),.co(c1_34_9)
);
wire c1_34_10, s1_34_10;
half_adder ha1_34_10 (
.a(A[30] & B[4]),.b(A[31] & B[3]),.p(s1_34_10),.g(c1_34_10)
);
wire c1_35_1, s1_35_1;
full_adder fa1_35_1 (
.a(A[4] & B[31]),.b(A[5] & B[30]),.c(A[6] & B[29]),.s(s1_35_1),.co(c1_35_1)
);
wire c1_35_2, s1_35_2;
full_adder fa1_35_2 (
.a(A[7] & B[28]),.b(A[8] & B[27]),.c(A[9] & B[26]),.s(s1_35_2),.co(c1_35_2)
);
wire c1_35_3, s1_35_3;
full_adder fa1_35_3 (
.a(A[10] & B[25]),.b(A[11] & B[24]),.c(A[12] & B[23]),.s(s1_35_3),.co(c1_35_3)
);
wire c1_35_4, s1_35_4;
full_adder fa1_35_4 (
.a(A[13] & B[22]),.b(A[14] & B[21]),.c(A[15] & B[20]),.s(s1_35_4),.co(c1_35_4)
);
wire c1_35_5, s1_35_5;
full_adder fa1_35_5 (
.a(A[16] & B[19]),.b(A[17] & B[18]),.c(A[18] & B[17]),.s(s1_35_5),.co(c1_35_5)
);
wire c1_35_6, s1_35_6;
full_adder fa1_35_6 (
.a(A[19] & B[16]),.b(A[20] & B[15]),.c(A[21] & B[14]),.s(s1_35_6),.co(c1_35_6)
);
wire c1_35_7, s1_35_7;
full_adder fa1_35_7 (
.a(A[22] & B[13]),.b(A[23] & B[12]),.c(A[24] & B[11]),.s(s1_35_7),.co(c1_35_7)
);
wire c1_35_8, s1_35_8;
full_adder fa1_35_8 (
.a(A[25] & B[10]),.b(A[26] & B[9]),.c(A[27] & B[8]),.s(s1_35_8),.co(c1_35_8)
);
wire c1_35_9, s1_35_9;
full_adder fa1_35_9 (
.a(A[28] & B[7]),.b(A[29] & B[6]),.c(A[30] & B[5]),.s(s1_35_9),.co(c1_35_9)
);
wire c1_36_1, s1_36_1;
full_adder fa1_36_1 (
.a(A[5] & B[31]),.b(A[6] & B[30]),.c(A[7] & B[29]),.s(s1_36_1),.co(c1_36_1)
);
wire c1_36_2, s1_36_2;
full_adder fa1_36_2 (
.a(A[8] & B[28]),.b(A[9] & B[27]),.c(A[10] & B[26]),.s(s1_36_2),.co(c1_36_2)
);
wire c1_36_3, s1_36_3;
full_adder fa1_36_3 (
.a(A[11] & B[25]),.b(A[12] & B[24]),.c(A[13] & B[23]),.s(s1_36_3),.co(c1_36_3)
);
wire c1_36_4, s1_36_4;
full_adder fa1_36_4 (
.a(A[14] & B[22]),.b(A[15] & B[21]),.c(A[16] & B[20]),.s(s1_36_4),.co(c1_36_4)
);
wire c1_36_5, s1_36_5;
full_adder fa1_36_5 (
.a(A[17] & B[19]),.b(A[18] & B[18]),.c(A[19] & B[17]),.s(s1_36_5),.co(c1_36_5)
);
wire c1_36_6, s1_36_6;
full_adder fa1_36_6 (
.a(A[20] & B[16]),.b(A[21] & B[15]),.c(A[22] & B[14]),.s(s1_36_6),.co(c1_36_6)
);
wire c1_36_7, s1_36_7;
full_adder fa1_36_7 (
.a(A[23] & B[13]),.b(A[24] & B[12]),.c(A[25] & B[11]),.s(s1_36_7),.co(c1_36_7)
);
wire c1_36_8, s1_36_8;
full_adder fa1_36_8 (
.a(A[26] & B[10]),.b(A[27] & B[9]),.c(A[28] & B[8]),.s(s1_36_8),.co(c1_36_8)
);
wire c1_36_9, s1_36_9;
full_adder fa1_36_9 (
.a(A[29] & B[7]),.b(A[30] & B[6]),.c(A[31] & B[5]),.s(s1_36_9),.co(c1_36_9)
);
wire c1_37_1, s1_37_1;
full_adder fa1_37_1 (
.a(A[6] & B[31]),.b(A[7] & B[30]),.c(A[8] & B[29]),.s(s1_37_1),.co(c1_37_1)
);
wire c1_37_2, s1_37_2;
full_adder fa1_37_2 (
.a(A[9] & B[28]),.b(A[10] & B[27]),.c(A[11] & B[26]),.s(s1_37_2),.co(c1_37_2)
);
wire c1_37_3, s1_37_3;
full_adder fa1_37_3 (
.a(A[12] & B[25]),.b(A[13] & B[24]),.c(A[14] & B[23]),.s(s1_37_3),.co(c1_37_3)
);
wire c1_37_4, s1_37_4;
full_adder fa1_37_4 (
.a(A[15] & B[22]),.b(A[16] & B[21]),.c(A[17] & B[20]),.s(s1_37_4),.co(c1_37_4)
);
wire c1_37_5, s1_37_5;
full_adder fa1_37_5 (
.a(A[18] & B[19]),.b(A[19] & B[18]),.c(A[20] & B[17]),.s(s1_37_5),.co(c1_37_5)
);
wire c1_37_6, s1_37_6;
full_adder fa1_37_6 (
.a(A[21] & B[16]),.b(A[22] & B[15]),.c(A[23] & B[14]),.s(s1_37_6),.co(c1_37_6)
);
wire c1_37_7, s1_37_7;
full_adder fa1_37_7 (
.a(A[24] & B[13]),.b(A[25] & B[12]),.c(A[26] & B[11]),.s(s1_37_7),.co(c1_37_7)
);
wire c1_37_8, s1_37_8;
full_adder fa1_37_8 (
.a(A[27] & B[10]),.b(A[28] & B[9]),.c(A[29] & B[8]),.s(s1_37_8),.co(c1_37_8)
);
wire c1_37_9, s1_37_9;
half_adder ha1_37_9 (
.a(A[30] & B[7]),.b(A[31] & B[6]),.p(s1_37_9),.g(c1_37_9)
);
wire c1_38_1, s1_38_1;
full_adder fa1_38_1 (
.a(A[7] & B[31]),.b(A[8] & B[30]),.c(A[9] & B[29]),.s(s1_38_1),.co(c1_38_1)
);
wire c1_38_2, s1_38_2;
full_adder fa1_38_2 (
.a(A[10] & B[28]),.b(A[11] & B[27]),.c(A[12] & B[26]),.s(s1_38_2),.co(c1_38_2)
);
wire c1_38_3, s1_38_3;
full_adder fa1_38_3 (
.a(A[13] & B[25]),.b(A[14] & B[24]),.c(A[15] & B[23]),.s(s1_38_3),.co(c1_38_3)
);
wire c1_38_4, s1_38_4;
full_adder fa1_38_4 (
.a(A[16] & B[22]),.b(A[17] & B[21]),.c(A[18] & B[20]),.s(s1_38_4),.co(c1_38_4)
);
wire c1_38_5, s1_38_5;
full_adder fa1_38_5 (
.a(A[19] & B[19]),.b(A[20] & B[18]),.c(A[21] & B[17]),.s(s1_38_5),.co(c1_38_5)
);
wire c1_38_6, s1_38_6;
full_adder fa1_38_6 (
.a(A[22] & B[16]),.b(A[23] & B[15]),.c(A[24] & B[14]),.s(s1_38_6),.co(c1_38_6)
);
wire c1_38_7, s1_38_7;
full_adder fa1_38_7 (
.a(A[25] & B[13]),.b(A[26] & B[12]),.c(A[27] & B[11]),.s(s1_38_7),.co(c1_38_7)
);
wire c1_38_8, s1_38_8;
full_adder fa1_38_8 (
.a(A[28] & B[10]),.b(A[29] & B[9]),.c(A[30] & B[8]),.s(s1_38_8),.co(c1_38_8)
);
wire c1_39_1, s1_39_1;
full_adder fa1_39_1 (
.a(A[8] & B[31]),.b(A[9] & B[30]),.c(A[10] & B[29]),.s(s1_39_1),.co(c1_39_1)
);
wire c1_39_2, s1_39_2;
full_adder fa1_39_2 (
.a(A[11] & B[28]),.b(A[12] & B[27]),.c(A[13] & B[26]),.s(s1_39_2),.co(c1_39_2)
);
wire c1_39_3, s1_39_3;
full_adder fa1_39_3 (
.a(A[14] & B[25]),.b(A[15] & B[24]),.c(A[16] & B[23]),.s(s1_39_3),.co(c1_39_3)
);
wire c1_39_4, s1_39_4;
full_adder fa1_39_4 (
.a(A[17] & B[22]),.b(A[18] & B[21]),.c(A[19] & B[20]),.s(s1_39_4),.co(c1_39_4)
);
wire c1_39_5, s1_39_5;
full_adder fa1_39_5 (
.a(A[20] & B[19]),.b(A[21] & B[18]),.c(A[22] & B[17]),.s(s1_39_5),.co(c1_39_5)
);
wire c1_39_6, s1_39_6;
full_adder fa1_39_6 (
.a(A[23] & B[16]),.b(A[24] & B[15]),.c(A[25] & B[14]),.s(s1_39_6),.co(c1_39_6)
);
wire c1_39_7, s1_39_7;
full_adder fa1_39_7 (
.a(A[26] & B[13]),.b(A[27] & B[12]),.c(A[28] & B[11]),.s(s1_39_7),.co(c1_39_7)
);
wire c1_39_8, s1_39_8;
full_adder fa1_39_8 (
.a(A[29] & B[10]),.b(A[30] & B[9]),.c(A[31] & B[8]),.s(s1_39_8),.co(c1_39_8)
);
wire c1_40_1, s1_40_1;
full_adder fa1_40_1 (
.a(A[9] & B[31]),.b(A[10] & B[30]),.c(A[11] & B[29]),.s(s1_40_1),.co(c1_40_1)
);
wire c1_40_2, s1_40_2;
full_adder fa1_40_2 (
.a(A[12] & B[28]),.b(A[13] & B[27]),.c(A[14] & B[26]),.s(s1_40_2),.co(c1_40_2)
);
wire c1_40_3, s1_40_3;
full_adder fa1_40_3 (
.a(A[15] & B[25]),.b(A[16] & B[24]),.c(A[17] & B[23]),.s(s1_40_3),.co(c1_40_3)
);
wire c1_40_4, s1_40_4;
full_adder fa1_40_4 (
.a(A[18] & B[22]),.b(A[19] & B[21]),.c(A[20] & B[20]),.s(s1_40_4),.co(c1_40_4)
);
wire c1_40_5, s1_40_5;
full_adder fa1_40_5 (
.a(A[21] & B[19]),.b(A[22] & B[18]),.c(A[23] & B[17]),.s(s1_40_5),.co(c1_40_5)
);
wire c1_40_6, s1_40_6;
full_adder fa1_40_6 (
.a(A[24] & B[16]),.b(A[25] & B[15]),.c(A[26] & B[14]),.s(s1_40_6),.co(c1_40_6)
);
wire c1_40_7, s1_40_7;
full_adder fa1_40_7 (
.a(A[27] & B[13]),.b(A[28] & B[12]),.c(A[29] & B[11]),.s(s1_40_7),.co(c1_40_7)
);
wire c1_40_8, s1_40_8;
half_adder ha1_40_8 (
.a(A[30] & B[10]),.b(A[31] & B[9]),.p(s1_40_8),.g(c1_40_8)
);
wire c1_41_1, s1_41_1;
full_adder fa1_41_1 (
.a(A[10] & B[31]),.b(A[11] & B[30]),.c(A[12] & B[29]),.s(s1_41_1),.co(c1_41_1)
);
wire c1_41_2, s1_41_2;
full_adder fa1_41_2 (
.a(A[13] & B[28]),.b(A[14] & B[27]),.c(A[15] & B[26]),.s(s1_41_2),.co(c1_41_2)
);
wire c1_41_3, s1_41_3;
full_adder fa1_41_3 (
.a(A[16] & B[25]),.b(A[17] & B[24]),.c(A[18] & B[23]),.s(s1_41_3),.co(c1_41_3)
);
wire c1_41_4, s1_41_4;
full_adder fa1_41_4 (
.a(A[19] & B[22]),.b(A[20] & B[21]),.c(A[21] & B[20]),.s(s1_41_4),.co(c1_41_4)
);
wire c1_41_5, s1_41_5;
full_adder fa1_41_5 (
.a(A[22] & B[19]),.b(A[23] & B[18]),.c(A[24] & B[17]),.s(s1_41_5),.co(c1_41_5)
);
wire c1_41_6, s1_41_6;
full_adder fa1_41_6 (
.a(A[25] & B[16]),.b(A[26] & B[15]),.c(A[27] & B[14]),.s(s1_41_6),.co(c1_41_6)
);
wire c1_41_7, s1_41_7;
full_adder fa1_41_7 (
.a(A[28] & B[13]),.b(A[29] & B[12]),.c(A[30] & B[11]),.s(s1_41_7),.co(c1_41_7)
);
wire c1_42_1, s1_42_1;
full_adder fa1_42_1 (
.a(A[11] & B[31]),.b(A[12] & B[30]),.c(A[13] & B[29]),.s(s1_42_1),.co(c1_42_1)
);
wire c1_42_2, s1_42_2;
full_adder fa1_42_2 (
.a(A[14] & B[28]),.b(A[15] & B[27]),.c(A[16] & B[26]),.s(s1_42_2),.co(c1_42_2)
);
wire c1_42_3, s1_42_3;
full_adder fa1_42_3 (
.a(A[17] & B[25]),.b(A[18] & B[24]),.c(A[19] & B[23]),.s(s1_42_3),.co(c1_42_3)
);
wire c1_42_4, s1_42_4;
full_adder fa1_42_4 (
.a(A[20] & B[22]),.b(A[21] & B[21]),.c(A[22] & B[20]),.s(s1_42_4),.co(c1_42_4)
);
wire c1_42_5, s1_42_5;
full_adder fa1_42_5 (
.a(A[23] & B[19]),.b(A[24] & B[18]),.c(A[25] & B[17]),.s(s1_42_5),.co(c1_42_5)
);
wire c1_42_6, s1_42_6;
full_adder fa1_42_6 (
.a(A[26] & B[16]),.b(A[27] & B[15]),.c(A[28] & B[14]),.s(s1_42_6),.co(c1_42_6)
);
wire c1_42_7, s1_42_7;
full_adder fa1_42_7 (
.a(A[29] & B[13]),.b(A[30] & B[12]),.c(A[31] & B[11]),.s(s1_42_7),.co(c1_42_7)
);
wire c1_43_1, s1_43_1;
full_adder fa1_43_1 (
.a(A[12] & B[31]),.b(A[13] & B[30]),.c(A[14] & B[29]),.s(s1_43_1),.co(c1_43_1)
);
wire c1_43_2, s1_43_2;
full_adder fa1_43_2 (
.a(A[15] & B[28]),.b(A[16] & B[27]),.c(A[17] & B[26]),.s(s1_43_2),.co(c1_43_2)
);
wire c1_43_3, s1_43_3;
full_adder fa1_43_3 (
.a(A[18] & B[25]),.b(A[19] & B[24]),.c(A[20] & B[23]),.s(s1_43_3),.co(c1_43_3)
);
wire c1_43_4, s1_43_4;
full_adder fa1_43_4 (
.a(A[21] & B[22]),.b(A[22] & B[21]),.c(A[23] & B[20]),.s(s1_43_4),.co(c1_43_4)
);
wire c1_43_5, s1_43_5;
full_adder fa1_43_5 (
.a(A[24] & B[19]),.b(A[25] & B[18]),.c(A[26] & B[17]),.s(s1_43_5),.co(c1_43_5)
);
wire c1_43_6, s1_43_6;
full_adder fa1_43_6 (
.a(A[27] & B[16]),.b(A[28] & B[15]),.c(A[29] & B[14]),.s(s1_43_6),.co(c1_43_6)
);
wire c1_43_7, s1_43_7;
half_adder ha1_43_7 (
.a(A[30] & B[13]),.b(A[31] & B[12]),.p(s1_43_7),.g(c1_43_7)
);
wire c1_44_1, s1_44_1;
full_adder fa1_44_1 (
.a(A[13] & B[31]),.b(A[14] & B[30]),.c(A[15] & B[29]),.s(s1_44_1),.co(c1_44_1)
);
wire c1_44_2, s1_44_2;
full_adder fa1_44_2 (
.a(A[16] & B[28]),.b(A[17] & B[27]),.c(A[18] & B[26]),.s(s1_44_2),.co(c1_44_2)
);
wire c1_44_3, s1_44_3;
full_adder fa1_44_3 (
.a(A[19] & B[25]),.b(A[20] & B[24]),.c(A[21] & B[23]),.s(s1_44_3),.co(c1_44_3)
);
wire c1_44_4, s1_44_4;
full_adder fa1_44_4 (
.a(A[22] & B[22]),.b(A[23] & B[21]),.c(A[24] & B[20]),.s(s1_44_4),.co(c1_44_4)
);
wire c1_44_5, s1_44_5;
full_adder fa1_44_5 (
.a(A[25] & B[19]),.b(A[26] & B[18]),.c(A[27] & B[17]),.s(s1_44_5),.co(c1_44_5)
);
wire c1_44_6, s1_44_6;
full_adder fa1_44_6 (
.a(A[28] & B[16]),.b(A[29] & B[15]),.c(A[30] & B[14]),.s(s1_44_6),.co(c1_44_6)
);
wire c1_45_1, s1_45_1;
full_adder fa1_45_1 (
.a(A[14] & B[31]),.b(A[15] & B[30]),.c(A[16] & B[29]),.s(s1_45_1),.co(c1_45_1)
);
wire c1_45_2, s1_45_2;
full_adder fa1_45_2 (
.a(A[17] & B[28]),.b(A[18] & B[27]),.c(A[19] & B[26]),.s(s1_45_2),.co(c1_45_2)
);
wire c1_45_3, s1_45_3;
full_adder fa1_45_3 (
.a(A[20] & B[25]),.b(A[21] & B[24]),.c(A[22] & B[23]),.s(s1_45_3),.co(c1_45_3)
);
wire c1_45_4, s1_45_4;
full_adder fa1_45_4 (
.a(A[23] & B[22]),.b(A[24] & B[21]),.c(A[25] & B[20]),.s(s1_45_4),.co(c1_45_4)
);
wire c1_45_5, s1_45_5;
full_adder fa1_45_5 (
.a(A[26] & B[19]),.b(A[27] & B[18]),.c(A[28] & B[17]),.s(s1_45_5),.co(c1_45_5)
);
wire c1_45_6, s1_45_6;
full_adder fa1_45_6 (
.a(A[29] & B[16]),.b(A[30] & B[15]),.c(A[31] & B[14]),.s(s1_45_6),.co(c1_45_6)
);
wire c1_46_1, s1_46_1;
full_adder fa1_46_1 (
.a(A[15] & B[31]),.b(A[16] & B[30]),.c(A[17] & B[29]),.s(s1_46_1),.co(c1_46_1)
);
wire c1_46_2, s1_46_2;
full_adder fa1_46_2 (
.a(A[18] & B[28]),.b(A[19] & B[27]),.c(A[20] & B[26]),.s(s1_46_2),.co(c1_46_2)
);
wire c1_46_3, s1_46_3;
full_adder fa1_46_3 (
.a(A[21] & B[25]),.b(A[22] & B[24]),.c(A[23] & B[23]),.s(s1_46_3),.co(c1_46_3)
);
wire c1_46_4, s1_46_4;
full_adder fa1_46_4 (
.a(A[24] & B[22]),.b(A[25] & B[21]),.c(A[26] & B[20]),.s(s1_46_4),.co(c1_46_4)
);
wire c1_46_5, s1_46_5;
full_adder fa1_46_5 (
.a(A[27] & B[19]),.b(A[28] & B[18]),.c(A[29] & B[17]),.s(s1_46_5),.co(c1_46_5)
);
wire c1_46_6, s1_46_6;
half_adder ha1_46_6 (
.a(A[30] & B[16]),.b(A[31] & B[15]),.p(s1_46_6),.g(c1_46_6)
);
wire c1_47_1, s1_47_1;
full_adder fa1_47_1 (
.a(A[16] & B[31]),.b(A[17] & B[30]),.c(A[18] & B[29]),.s(s1_47_1),.co(c1_47_1)
);
wire c1_47_2, s1_47_2;
full_adder fa1_47_2 (
.a(A[19] & B[28]),.b(A[20] & B[27]),.c(A[21] & B[26]),.s(s1_47_2),.co(c1_47_2)
);
wire c1_47_3, s1_47_3;
full_adder fa1_47_3 (
.a(A[22] & B[25]),.b(A[23] & B[24]),.c(A[24] & B[23]),.s(s1_47_3),.co(c1_47_3)
);
wire c1_47_4, s1_47_4;
full_adder fa1_47_4 (
.a(A[25] & B[22]),.b(A[26] & B[21]),.c(A[27] & B[20]),.s(s1_47_4),.co(c1_47_4)
);
wire c1_47_5, s1_47_5;
full_adder fa1_47_5 (
.a(A[28] & B[19]),.b(A[29] & B[18]),.c(A[30] & B[17]),.s(s1_47_5),.co(c1_47_5)
);
wire c1_48_1, s1_48_1;
full_adder fa1_48_1 (
.a(A[17] & B[31]),.b(A[18] & B[30]),.c(A[19] & B[29]),.s(s1_48_1),.co(c1_48_1)
);
wire c1_48_2, s1_48_2;
full_adder fa1_48_2 (
.a(A[20] & B[28]),.b(A[21] & B[27]),.c(A[22] & B[26]),.s(s1_48_2),.co(c1_48_2)
);
wire c1_48_3, s1_48_3;
full_adder fa1_48_3 (
.a(A[23] & B[25]),.b(A[24] & B[24]),.c(A[25] & B[23]),.s(s1_48_3),.co(c1_48_3)
);
wire c1_48_4, s1_48_4;
full_adder fa1_48_4 (
.a(A[26] & B[22]),.b(A[27] & B[21]),.c(A[28] & B[20]),.s(s1_48_4),.co(c1_48_4)
);
wire c1_48_5, s1_48_5;
full_adder fa1_48_5 (
.a(A[29] & B[19]),.b(A[30] & B[18]),.c(A[31] & B[17]),.s(s1_48_5),.co(c1_48_5)
);
wire c1_49_1, s1_49_1;
full_adder fa1_49_1 (
.a(A[18] & B[31]),.b(A[19] & B[30]),.c(A[20] & B[29]),.s(s1_49_1),.co(c1_49_1)
);
wire c1_49_2, s1_49_2;
full_adder fa1_49_2 (
.a(A[21] & B[28]),.b(A[22] & B[27]),.c(A[23] & B[26]),.s(s1_49_2),.co(c1_49_2)
);
wire c1_49_3, s1_49_3;
full_adder fa1_49_3 (
.a(A[24] & B[25]),.b(A[25] & B[24]),.c(A[26] & B[23]),.s(s1_49_3),.co(c1_49_3)
);
wire c1_49_4, s1_49_4;
full_adder fa1_49_4 (
.a(A[27] & B[22]),.b(A[28] & B[21]),.c(A[29] & B[20]),.s(s1_49_4),.co(c1_49_4)
);
wire c1_49_5, s1_49_5;
half_adder ha1_49_5 (
.a(A[30] & B[19]),.b(A[31] & B[18]),.p(s1_49_5),.g(c1_49_5)
);
wire c1_50_1, s1_50_1;
full_adder fa1_50_1 (
.a(A[19] & B[31]),.b(A[20] & B[30]),.c(A[21] & B[29]),.s(s1_50_1),.co(c1_50_1)
);
wire c1_50_2, s1_50_2;
full_adder fa1_50_2 (
.a(A[22] & B[28]),.b(A[23] & B[27]),.c(A[24] & B[26]),.s(s1_50_2),.co(c1_50_2)
);
wire c1_50_3, s1_50_3;
full_adder fa1_50_3 (
.a(A[25] & B[25]),.b(A[26] & B[24]),.c(A[27] & B[23]),.s(s1_50_3),.co(c1_50_3)
);
wire c1_50_4, s1_50_4;
full_adder fa1_50_4 (
.a(A[28] & B[22]),.b(A[29] & B[21]),.c(A[30] & B[20]),.s(s1_50_4),.co(c1_50_4)
);
wire c1_51_1, s1_51_1;
full_adder fa1_51_1 (
.a(A[20] & B[31]),.b(A[21] & B[30]),.c(A[22] & B[29]),.s(s1_51_1),.co(c1_51_1)
);
wire c1_51_2, s1_51_2;
full_adder fa1_51_2 (
.a(A[23] & B[28]),.b(A[24] & B[27]),.c(A[25] & B[26]),.s(s1_51_2),.co(c1_51_2)
);
wire c1_51_3, s1_51_3;
full_adder fa1_51_3 (
.a(A[26] & B[25]),.b(A[27] & B[24]),.c(A[28] & B[23]),.s(s1_51_3),.co(c1_51_3)
);
wire c1_51_4, s1_51_4;
full_adder fa1_51_4 (
.a(A[29] & B[22]),.b(A[30] & B[21]),.c(A[31] & B[20]),.s(s1_51_4),.co(c1_51_4)
);
wire c1_52_1, s1_52_1;
full_adder fa1_52_1 (
.a(A[21] & B[31]),.b(A[22] & B[30]),.c(A[23] & B[29]),.s(s1_52_1),.co(c1_52_1)
);
wire c1_52_2, s1_52_2;
full_adder fa1_52_2 (
.a(A[24] & B[28]),.b(A[25] & B[27]),.c(A[26] & B[26]),.s(s1_52_2),.co(c1_52_2)
);
wire c1_52_3, s1_52_3;
full_adder fa1_52_3 (
.a(A[27] & B[25]),.b(A[28] & B[24]),.c(A[29] & B[23]),.s(s1_52_3),.co(c1_52_3)
);
wire c1_52_4, s1_52_4;
half_adder ha1_52_4 (
.a(A[30] & B[22]),.b(A[31] & B[21]),.p(s1_52_4),.g(c1_52_4)
);
wire c1_53_1, s1_53_1;
full_adder fa1_53_1 (
.a(A[22] & B[31]),.b(A[23] & B[30]),.c(A[24] & B[29]),.s(s1_53_1),.co(c1_53_1)
);
wire c1_53_2, s1_53_2;
full_adder fa1_53_2 (
.a(A[25] & B[28]),.b(A[26] & B[27]),.c(A[27] & B[26]),.s(s1_53_2),.co(c1_53_2)
);
wire c1_53_3, s1_53_3;
full_adder fa1_53_3 (
.a(A[28] & B[25]),.b(A[29] & B[24]),.c(A[30] & B[23]),.s(s1_53_3),.co(c1_53_3)
);
wire c1_54_1, s1_54_1;
full_adder fa1_54_1 (
.a(A[23] & B[31]),.b(A[24] & B[30]),.c(A[25] & B[29]),.s(s1_54_1),.co(c1_54_1)
);
wire c1_54_2, s1_54_2;
full_adder fa1_54_2 (
.a(A[26] & B[28]),.b(A[27] & B[27]),.c(A[28] & B[26]),.s(s1_54_2),.co(c1_54_2)
);
wire c1_54_3, s1_54_3;
full_adder fa1_54_3 (
.a(A[29] & B[25]),.b(A[30] & B[24]),.c(A[31] & B[23]),.s(s1_54_3),.co(c1_54_3)
);
wire c1_55_1, s1_55_1;
full_adder fa1_55_1 (
.a(A[24] & B[31]),.b(A[25] & B[30]),.c(A[26] & B[29]),.s(s1_55_1),.co(c1_55_1)
);
wire c1_55_2, s1_55_2;
full_adder fa1_55_2 (
.a(A[27] & B[28]),.b(A[28] & B[27]),.c(A[29] & B[26]),.s(s1_55_2),.co(c1_55_2)
);
wire c1_55_3, s1_55_3;
half_adder ha1_55_3 (
.a(A[30] & B[25]),.b(A[31] & B[24]),.p(s1_55_3),.g(c1_55_3)
);
wire c1_56_1, s1_56_1;
full_adder fa1_56_1 (
.a(A[25] & B[31]),.b(A[26] & B[30]),.c(A[27] & B[29]),.s(s1_56_1),.co(c1_56_1)
);
wire c1_56_2, s1_56_2;
full_adder fa1_56_2 (
.a(A[28] & B[28]),.b(A[29] & B[27]),.c(A[30] & B[26]),.s(s1_56_2),.co(c1_56_2)
);
wire c1_57_1, s1_57_1;
full_adder fa1_57_1 (
.a(A[26] & B[31]),.b(A[27] & B[30]),.c(A[28] & B[29]),.s(s1_57_1),.co(c1_57_1)
);
wire c1_57_2, s1_57_2;
full_adder fa1_57_2 (
.a(A[29] & B[28]),.b(A[30] & B[27]),.c(A[31] & B[26]),.s(s1_57_2),.co(c1_57_2)
);
wire c1_58_1, s1_58_1;
full_adder fa1_58_1 (
.a(A[27] & B[31]),.b(A[28] & B[30]),.c(A[29] & B[29]),.s(s1_58_1),.co(c1_58_1)
);
wire c1_58_2, s1_58_2;
half_adder ha1_58_2 (
.a(A[30] & B[28]),.b(A[31] & B[27]),.p(s1_58_2),.g(c1_58_2)
);
wire c1_59_1, s1_59_1;
full_adder fa1_59_1 (
.a(A[28] & B[31]),.b(A[29] & B[30]),.c(A[30] & B[29]),.s(s1_59_1),.co(c1_59_1)
);
wire c1_60_1, s1_60_1;
full_adder fa1_60_1 (
.a(A[29] & B[31]),.b(A[30] & B[30]),.c(A[31] & B[29]),.s(s1_60_1),.co(c1_60_1)
);
wire c1_61_1, s1_61_1;
half_adder ha1_61_1 (
.a(A[30] & B[31]),.b(A[31] & B[30]),.p(s1_61_1),.g(c1_61_1)
);
wire c2_2_1, s2_2_1;
half_adder ha2_2_1 (
.a(s1_2_1),.b(c1_1_1),.p(s2_2_1),.g(c2_2_1)
);
wire c2_3_1, s2_3_1;
full_adder fa2_3_1 (
.a(A[3] & B[0]),.b(s1_3_1),.c(c1_2_1),.s(s2_3_1),.co(c2_3_1)
);
wire c2_4_1, s2_4_1;
full_adder fa2_4_1 (
.a(s1_4_2),.b(s1_4_1),.c(c1_3_1),.s(s2_4_1),.co(c2_4_1)
);
wire c2_5_1, s2_5_1;
full_adder fa2_5_1 (
.a(s1_5_2),.b(s1_5_1),.c(c1_4_2),.s(s2_5_1),.co(c2_5_1)
);
wire c2_6_1, s2_6_1;
full_adder fa2_6_1 (
.a(A[6] & B[0]),.b(s1_6_2),.c(s1_6_1),.s(s2_6_1),.co(c2_6_1)
);
wire c2_6_2, s2_6_2;
half_adder ha2_6_2 (
.a(c1_5_2),.b(c1_5_1),.p(s2_6_2),.g(c2_6_2)
);
wire c2_7_1, s2_7_1;
full_adder fa2_7_1 (
.a(s1_7_3),.b(s1_7_2),.c(s1_7_1),.s(s2_7_1),.co(c2_7_1)
);
wire c2_7_2, s2_7_2;
half_adder ha2_7_2 (
.a(c1_6_2),.b(c1_6_1),.p(s2_7_2),.g(c2_7_2)
);
wire c2_8_1, s2_8_1;
full_adder fa2_8_1 (
.a(s1_8_3),.b(s1_8_2),.c(s1_8_1),.s(s2_8_1),.co(c2_8_1)
);
wire c2_8_2, s2_8_2;
full_adder fa2_8_2 (
.a(c1_7_3),.b(c1_7_2),.c(c1_7_1),.s(s2_8_2),.co(c2_8_2)
);
wire c2_9_1, s2_9_1;
full_adder fa2_9_1 (
.a(A[9] & B[0]),.b(s1_9_3),.c(s1_9_2),.s(s2_9_1),.co(c2_9_1)
);
wire c2_9_2, s2_9_2;
full_adder fa2_9_2 (
.a(s1_9_1),.b(c1_8_3),.c(c1_8_2),.s(s2_9_2),.co(c2_9_2)
);
wire c2_10_1, s2_10_1;
full_adder fa2_10_1 (
.a(s1_10_4),.b(s1_10_3),.c(s1_10_2),.s(s2_10_1),.co(c2_10_1)
);
wire c2_10_2, s2_10_2;
full_adder fa2_10_2 (
.a(s1_10_1),.b(c1_9_3),.c(c1_9_2),.s(s2_10_2),.co(c2_10_2)
);
wire c2_11_1, s2_11_1;
full_adder fa2_11_1 (
.a(s1_11_4),.b(s1_11_3),.c(s1_11_2),.s(s2_11_1),.co(c2_11_1)
);
wire c2_11_2, s2_11_2;
full_adder fa2_11_2 (
.a(s1_11_1),.b(c1_10_4),.c(c1_10_3),.s(s2_11_2),.co(c2_11_2)
);
wire c2_11_3, s2_11_3;
half_adder ha2_11_3 (
.a(c1_10_2),.b(c1_10_1),.p(s2_11_3),.g(c2_11_3)
);
wire c2_12_1, s2_12_1;
full_adder fa2_12_1 (
.a(A[12] & B[0]),.b(s1_12_4),.c(s1_12_3),.s(s2_12_1),.co(c2_12_1)
);
wire c2_12_2, s2_12_2;
full_adder fa2_12_2 (
.a(s1_12_2),.b(s1_12_1),.c(c1_11_4),.s(s2_12_2),.co(c2_12_2)
);
wire c2_12_3, s2_12_3;
full_adder fa2_12_3 (
.a(c1_11_3),.b(c1_11_2),.c(c1_11_1),.s(s2_12_3),.co(c2_12_3)
);
wire c2_13_1, s2_13_1;
full_adder fa2_13_1 (
.a(s1_13_5),.b(s1_13_4),.c(s1_13_3),.s(s2_13_1),.co(c2_13_1)
);
wire c2_13_2, s2_13_2;
full_adder fa2_13_2 (
.a(s1_13_2),.b(s1_13_1),.c(c1_12_4),.s(s2_13_2),.co(c2_13_2)
);
wire c2_13_3, s2_13_3;
full_adder fa2_13_3 (
.a(c1_12_3),.b(c1_12_2),.c(c1_12_1),.s(s2_13_3),.co(c2_13_3)
);
wire c2_14_1, s2_14_1;
full_adder fa2_14_1 (
.a(s1_14_5),.b(s1_14_4),.c(s1_14_3),.s(s2_14_1),.co(c2_14_1)
);
wire c2_14_2, s2_14_2;
full_adder fa2_14_2 (
.a(s1_14_2),.b(s1_14_1),.c(c1_13_5),.s(s2_14_2),.co(c2_14_2)
);
wire c2_14_3, s2_14_3;
full_adder fa2_14_3 (
.a(c1_13_4),.b(c1_13_3),.c(c1_13_2),.s(s2_14_3),.co(c2_14_3)
);
wire c2_15_1, s2_15_1;
full_adder fa2_15_1 (
.a(A[15] & B[0]),.b(s1_15_5),.c(s1_15_4),.s(s2_15_1),.co(c2_15_1)
);
wire c2_15_2, s2_15_2;
full_adder fa2_15_2 (
.a(s1_15_3),.b(s1_15_2),.c(s1_15_1),.s(s2_15_2),.co(c2_15_2)
);
wire c2_15_3, s2_15_3;
full_adder fa2_15_3 (
.a(c1_14_5),.b(c1_14_4),.c(c1_14_3),.s(s2_15_3),.co(c2_15_3)
);
wire c2_15_4, s2_15_4;
half_adder ha2_15_4 (
.a(c1_14_2),.b(c1_14_1),.p(s2_15_4),.g(c2_15_4)
);
wire c2_16_1, s2_16_1;
full_adder fa2_16_1 (
.a(s1_16_6),.b(s1_16_5),.c(s1_16_4),.s(s2_16_1),.co(c2_16_1)
);
wire c2_16_2, s2_16_2;
full_adder fa2_16_2 (
.a(s1_16_3),.b(s1_16_2),.c(s1_16_1),.s(s2_16_2),.co(c2_16_2)
);
wire c2_16_3, s2_16_3;
full_adder fa2_16_3 (
.a(c1_15_5),.b(c1_15_4),.c(c1_15_3),.s(s2_16_3),.co(c2_16_3)
);
wire c2_16_4, s2_16_4;
half_adder ha2_16_4 (
.a(c1_15_2),.b(c1_15_1),.p(s2_16_4),.g(c2_16_4)
);
wire c2_17_1, s2_17_1;
full_adder fa2_17_1 (
.a(s1_17_6),.b(s1_17_5),.c(s1_17_4),.s(s2_17_1),.co(c2_17_1)
);
wire c2_17_2, s2_17_2;
full_adder fa2_17_2 (
.a(s1_17_3),.b(s1_17_2),.c(s1_17_1),.s(s2_17_2),.co(c2_17_2)
);
wire c2_17_3, s2_17_3;
full_adder fa2_17_3 (
.a(c1_16_6),.b(c1_16_5),.c(c1_16_4),.s(s2_17_3),.co(c2_17_3)
);
wire c2_17_4, s2_17_4;
full_adder fa2_17_4 (
.a(c1_16_3),.b(c1_16_2),.c(c1_16_1),.s(s2_17_4),.co(c2_17_4)
);
wire c2_18_1, s2_18_1;
full_adder fa2_18_1 (
.a(A[18] & B[0]),.b(s1_18_6),.c(s1_18_5),.s(s2_18_1),.co(c2_18_1)
);
wire c2_18_2, s2_18_2;
full_adder fa2_18_2 (
.a(s1_18_4),.b(s1_18_3),.c(s1_18_2),.s(s2_18_2),.co(c2_18_2)
);
wire c2_18_3, s2_18_3;
full_adder fa2_18_3 (
.a(s1_18_1),.b(c1_17_6),.c(c1_17_5),.s(s2_18_3),.co(c2_18_3)
);
wire c2_18_4, s2_18_4;
full_adder fa2_18_4 (
.a(c1_17_4),.b(c1_17_3),.c(c1_17_2),.s(s2_18_4),.co(c2_18_4)
);
wire c2_19_1, s2_19_1;
full_adder fa2_19_1 (
.a(s1_19_7),.b(s1_19_6),.c(s1_19_5),.s(s2_19_1),.co(c2_19_1)
);
wire c2_19_2, s2_19_2;
full_adder fa2_19_2 (
.a(s1_19_4),.b(s1_19_3),.c(s1_19_2),.s(s2_19_2),.co(c2_19_2)
);
wire c2_19_3, s2_19_3;
full_adder fa2_19_3 (
.a(s1_19_1),.b(c1_18_6),.c(c1_18_5),.s(s2_19_3),.co(c2_19_3)
);
wire c2_19_4, s2_19_4;
full_adder fa2_19_4 (
.a(c1_18_4),.b(c1_18_3),.c(c1_18_2),.s(s2_19_4),.co(c2_19_4)
);
wire c2_20_1, s2_20_1;
full_adder fa2_20_1 (
.a(s1_20_7),.b(s1_20_6),.c(s1_20_5),.s(s2_20_1),.co(c2_20_1)
);
wire c2_20_2, s2_20_2;
full_adder fa2_20_2 (
.a(s1_20_4),.b(s1_20_3),.c(s1_20_2),.s(s2_20_2),.co(c2_20_2)
);
wire c2_20_3, s2_20_3;
full_adder fa2_20_3 (
.a(s1_20_1),.b(c1_19_7),.c(c1_19_6),.s(s2_20_3),.co(c2_20_3)
);
wire c2_20_4, s2_20_4;
full_adder fa2_20_4 (
.a(c1_19_5),.b(c1_19_4),.c(c1_19_3),.s(s2_20_4),.co(c2_20_4)
);
wire c2_20_5, s2_20_5;
half_adder ha2_20_5 (
.a(c1_19_2),.b(c1_19_1),.p(s2_20_5),.g(c2_20_5)
);
wire c2_21_1, s2_21_1;
full_adder fa2_21_1 (
.a(A[21] & B[0]),.b(s1_21_7),.c(s1_21_6),.s(s2_21_1),.co(c2_21_1)
);
wire c2_21_2, s2_21_2;
full_adder fa2_21_2 (
.a(s1_21_5),.b(s1_21_4),.c(s1_21_3),.s(s2_21_2),.co(c2_21_2)
);
wire c2_21_3, s2_21_3;
full_adder fa2_21_3 (
.a(s1_21_2),.b(s1_21_1),.c(c1_20_7),.s(s2_21_3),.co(c2_21_3)
);
wire c2_21_4, s2_21_4;
full_adder fa2_21_4 (
.a(c1_20_6),.b(c1_20_5),.c(c1_20_4),.s(s2_21_4),.co(c2_21_4)
);
wire c2_21_5, s2_21_5;
full_adder fa2_21_5 (
.a(c1_20_3),.b(c1_20_2),.c(c1_20_1),.s(s2_21_5),.co(c2_21_5)
);
wire c2_22_1, s2_22_1;
full_adder fa2_22_1 (
.a(s1_22_8),.b(s1_22_7),.c(s1_22_6),.s(s2_22_1),.co(c2_22_1)
);
wire c2_22_2, s2_22_2;
full_adder fa2_22_2 (
.a(s1_22_5),.b(s1_22_4),.c(s1_22_3),.s(s2_22_2),.co(c2_22_2)
);
wire c2_22_3, s2_22_3;
full_adder fa2_22_3 (
.a(s1_22_2),.b(s1_22_1),.c(c1_21_7),.s(s2_22_3),.co(c2_22_3)
);
wire c2_22_4, s2_22_4;
full_adder fa2_22_4 (
.a(c1_21_6),.b(c1_21_5),.c(c1_21_4),.s(s2_22_4),.co(c2_22_4)
);
wire c2_22_5, s2_22_5;
full_adder fa2_22_5 (
.a(c1_21_3),.b(c1_21_2),.c(c1_21_1),.s(s2_22_5),.co(c2_22_5)
);
wire c2_23_1, s2_23_1;
full_adder fa2_23_1 (
.a(s1_23_8),.b(s1_23_7),.c(s1_23_6),.s(s2_23_1),.co(c2_23_1)
);
wire c2_23_2, s2_23_2;
full_adder fa2_23_2 (
.a(s1_23_5),.b(s1_23_4),.c(s1_23_3),.s(s2_23_2),.co(c2_23_2)
);
wire c2_23_3, s2_23_3;
full_adder fa2_23_3 (
.a(s1_23_2),.b(s1_23_1),.c(c1_22_8),.s(s2_23_3),.co(c2_23_3)
);
wire c2_23_4, s2_23_4;
full_adder fa2_23_4 (
.a(c1_22_7),.b(c1_22_6),.c(c1_22_5),.s(s2_23_4),.co(c2_23_4)
);
wire c2_23_5, s2_23_5;
full_adder fa2_23_5 (
.a(c1_22_4),.b(c1_22_3),.c(c1_22_2),.s(s2_23_5),.co(c2_23_5)
);
wire c2_24_1, s2_24_1;
full_adder fa2_24_1 (
.a(A[24] & B[0]),.b(s1_24_8),.c(s1_24_7),.s(s2_24_1),.co(c2_24_1)
);
wire c2_24_2, s2_24_2;
full_adder fa2_24_2 (
.a(s1_24_6),.b(s1_24_5),.c(s1_24_4),.s(s2_24_2),.co(c2_24_2)
);
wire c2_24_3, s2_24_3;
full_adder fa2_24_3 (
.a(s1_24_3),.b(s1_24_2),.c(s1_24_1),.s(s2_24_3),.co(c2_24_3)
);
wire c2_24_4, s2_24_4;
full_adder fa2_24_4 (
.a(c1_23_8),.b(c1_23_7),.c(c1_23_6),.s(s2_24_4),.co(c2_24_4)
);
wire c2_24_5, s2_24_5;
full_adder fa2_24_5 (
.a(c1_23_5),.b(c1_23_4),.c(c1_23_3),.s(s2_24_5),.co(c2_24_5)
);
wire c2_24_6, s2_24_6;
half_adder ha2_24_6 (
.a(c1_23_2),.b(c1_23_1),.p(s2_24_6),.g(c2_24_6)
);
wire c2_25_1, s2_25_1;
full_adder fa2_25_1 (
.a(s1_25_9),.b(s1_25_8),.c(s1_25_7),.s(s2_25_1),.co(c2_25_1)
);
wire c2_25_2, s2_25_2;
full_adder fa2_25_2 (
.a(s1_25_6),.b(s1_25_5),.c(s1_25_4),.s(s2_25_2),.co(c2_25_2)
);
wire c2_25_3, s2_25_3;
full_adder fa2_25_3 (
.a(s1_25_3),.b(s1_25_2),.c(s1_25_1),.s(s2_25_3),.co(c2_25_3)
);
wire c2_25_4, s2_25_4;
full_adder fa2_25_4 (
.a(c1_24_8),.b(c1_24_7),.c(c1_24_6),.s(s2_25_4),.co(c2_25_4)
);
wire c2_25_5, s2_25_5;
full_adder fa2_25_5 (
.a(c1_24_5),.b(c1_24_4),.c(c1_24_3),.s(s2_25_5),.co(c2_25_5)
);
wire c2_25_6, s2_25_6;
half_adder ha2_25_6 (
.a(c1_24_2),.b(c1_24_1),.p(s2_25_6),.g(c2_25_6)
);
wire c2_26_1, s2_26_1;
full_adder fa2_26_1 (
.a(s1_26_9),.b(s1_26_8),.c(s1_26_7),.s(s2_26_1),.co(c2_26_1)
);
wire c2_26_2, s2_26_2;
full_adder fa2_26_2 (
.a(s1_26_6),.b(s1_26_5),.c(s1_26_4),.s(s2_26_2),.co(c2_26_2)
);
wire c2_26_3, s2_26_3;
full_adder fa2_26_3 (
.a(s1_26_3),.b(s1_26_2),.c(s1_26_1),.s(s2_26_3),.co(c2_26_3)
);
wire c2_26_4, s2_26_4;
full_adder fa2_26_4 (
.a(c1_25_9),.b(c1_25_8),.c(c1_25_7),.s(s2_26_4),.co(c2_26_4)
);
wire c2_26_5, s2_26_5;
full_adder fa2_26_5 (
.a(c1_25_6),.b(c1_25_5),.c(c1_25_4),.s(s2_26_5),.co(c2_26_5)
);
wire c2_26_6, s2_26_6;
full_adder fa2_26_6 (
.a(c1_25_3),.b(c1_25_2),.c(c1_25_1),.s(s2_26_6),.co(c2_26_6)
);
wire c2_27_1, s2_27_1;
full_adder fa2_27_1 (
.a(A[27] & B[0]),.b(s1_27_9),.c(s1_27_8),.s(s2_27_1),.co(c2_27_1)
);
wire c2_27_2, s2_27_2;
full_adder fa2_27_2 (
.a(s1_27_7),.b(s1_27_6),.c(s1_27_5),.s(s2_27_2),.co(c2_27_2)
);
wire c2_27_3, s2_27_3;
full_adder fa2_27_3 (
.a(s1_27_4),.b(s1_27_3),.c(s1_27_2),.s(s2_27_3),.co(c2_27_3)
);
wire c2_27_4, s2_27_4;
full_adder fa2_27_4 (
.a(s1_27_1),.b(c1_26_9),.c(c1_26_8),.s(s2_27_4),.co(c2_27_4)
);
wire c2_27_5, s2_27_5;
full_adder fa2_27_5 (
.a(c1_26_7),.b(c1_26_6),.c(c1_26_5),.s(s2_27_5),.co(c2_27_5)
);
wire c2_27_6, s2_27_6;
full_adder fa2_27_6 (
.a(c1_26_4),.b(c1_26_3),.c(c1_26_2),.s(s2_27_6),.co(c2_27_6)
);
wire c2_28_1, s2_28_1;
full_adder fa2_28_1 (
.a(s1_28_10),.b(s1_28_9),.c(s1_28_8),.s(s2_28_1),.co(c2_28_1)
);
wire c2_28_2, s2_28_2;
full_adder fa2_28_2 (
.a(s1_28_7),.b(s1_28_6),.c(s1_28_5),.s(s2_28_2),.co(c2_28_2)
);
wire c2_28_3, s2_28_3;
full_adder fa2_28_3 (
.a(s1_28_4),.b(s1_28_3),.c(s1_28_2),.s(s2_28_3),.co(c2_28_3)
);
wire c2_28_4, s2_28_4;
full_adder fa2_28_4 (
.a(s1_28_1),.b(c1_27_9),.c(c1_27_8),.s(s2_28_4),.co(c2_28_4)
);
wire c2_28_5, s2_28_5;
full_adder fa2_28_5 (
.a(c1_27_7),.b(c1_27_6),.c(c1_27_5),.s(s2_28_5),.co(c2_28_5)
);
wire c2_28_6, s2_28_6;
full_adder fa2_28_6 (
.a(c1_27_4),.b(c1_27_3),.c(c1_27_2),.s(s2_28_6),.co(c2_28_6)
);
wire c2_29_1, s2_29_1;
full_adder fa2_29_1 (
.a(s1_29_10),.b(s1_29_9),.c(s1_29_8),.s(s2_29_1),.co(c2_29_1)
);
wire c2_29_2, s2_29_2;
full_adder fa2_29_2 (
.a(s1_29_7),.b(s1_29_6),.c(s1_29_5),.s(s2_29_2),.co(c2_29_2)
);
wire c2_29_3, s2_29_3;
full_adder fa2_29_3 (
.a(s1_29_4),.b(s1_29_3),.c(s1_29_2),.s(s2_29_3),.co(c2_29_3)
);
wire c2_29_4, s2_29_4;
full_adder fa2_29_4 (
.a(s1_29_1),.b(c1_28_10),.c(c1_28_9),.s(s2_29_4),.co(c2_29_4)
);
wire c2_29_5, s2_29_5;
full_adder fa2_29_5 (
.a(c1_28_8),.b(c1_28_7),.c(c1_28_6),.s(s2_29_5),.co(c2_29_5)
);
wire c2_29_6, s2_29_6;
full_adder fa2_29_6 (
.a(c1_28_5),.b(c1_28_4),.c(c1_28_3),.s(s2_29_6),.co(c2_29_6)
);
wire c2_29_7, s2_29_7;
half_adder ha2_29_7 (
.a(c1_28_2),.b(c1_28_1),.p(s2_29_7),.g(c2_29_7)
);
wire c2_30_1, s2_30_1;
full_adder fa2_30_1 (
.a(A[30] & B[0]),.b(s1_30_10),.c(s1_30_9),.s(s2_30_1),.co(c2_30_1)
);
wire c2_30_2, s2_30_2;
full_adder fa2_30_2 (
.a(s1_30_8),.b(s1_30_7),.c(s1_30_6),.s(s2_30_2),.co(c2_30_2)
);
wire c2_30_3, s2_30_3;
full_adder fa2_30_3 (
.a(s1_30_5),.b(s1_30_4),.c(s1_30_3),.s(s2_30_3),.co(c2_30_3)
);
wire c2_30_4, s2_30_4;
full_adder fa2_30_4 (
.a(s1_30_2),.b(s1_30_1),.c(c1_29_10),.s(s2_30_4),.co(c2_30_4)
);
wire c2_30_5, s2_30_5;
full_adder fa2_30_5 (
.a(c1_29_9),.b(c1_29_8),.c(c1_29_7),.s(s2_30_5),.co(c2_30_5)
);
wire c2_30_6, s2_30_6;
full_adder fa2_30_6 (
.a(c1_29_6),.b(c1_29_5),.c(c1_29_4),.s(s2_30_6),.co(c2_30_6)
);
wire c2_30_7, s2_30_7;
full_adder fa2_30_7 (
.a(c1_29_3),.b(c1_29_2),.c(c1_29_1),.s(s2_30_7),.co(c2_30_7)
);
wire c2_31_1, s2_31_1;
full_adder fa2_31_1 (
.a(s1_31_11),.b(s1_31_10),.c(s1_31_9),.s(s2_31_1),.co(c2_31_1)
);
wire c2_31_2, s2_31_2;
full_adder fa2_31_2 (
.a(s1_31_8),.b(s1_31_7),.c(s1_31_6),.s(s2_31_2),.co(c2_31_2)
);
wire c2_31_3, s2_31_3;
full_adder fa2_31_3 (
.a(s1_31_5),.b(s1_31_4),.c(s1_31_3),.s(s2_31_3),.co(c2_31_3)
);
wire c2_31_4, s2_31_4;
full_adder fa2_31_4 (
.a(s1_31_2),.b(s1_31_1),.c(c1_30_10),.s(s2_31_4),.co(c2_31_4)
);
wire c2_31_5, s2_31_5;
full_adder fa2_31_5 (
.a(c1_30_9),.b(c1_30_8),.c(c1_30_7),.s(s2_31_5),.co(c2_31_5)
);
wire c2_31_6, s2_31_6;
full_adder fa2_31_6 (
.a(c1_30_6),.b(c1_30_5),.c(c1_30_4),.s(s2_31_6),.co(c2_31_6)
);
wire c2_31_7, s2_31_7;
full_adder fa2_31_7 (
.a(c1_30_3),.b(c1_30_2),.c(c1_30_1),.s(s2_31_7),.co(c2_31_7)
);
wire c2_32_1, s2_32_1;
full_adder fa2_32_1 (
.a(A[31] & B[1]),.b(s1_32_10),.c(s1_32_9),.s(s2_32_1),.co(c2_32_1)
);
wire c2_32_2, s2_32_2;
full_adder fa2_32_2 (
.a(s1_32_8),.b(s1_32_7),.c(s1_32_6),.s(s2_32_2),.co(c2_32_2)
);
wire c2_32_3, s2_32_3;
full_adder fa2_32_3 (
.a(s1_32_5),.b(s1_32_4),.c(s1_32_3),.s(s2_32_3),.co(c2_32_3)
);
wire c2_32_4, s2_32_4;
full_adder fa2_32_4 (
.a(s1_32_2),.b(s1_32_1),.c(c1_31_11),.s(s2_32_4),.co(c2_32_4)
);
wire c2_32_5, s2_32_5;
full_adder fa2_32_5 (
.a(c1_31_10),.b(c1_31_9),.c(c1_31_8),.s(s2_32_5),.co(c2_32_5)
);
wire c2_32_6, s2_32_6;
full_adder fa2_32_6 (
.a(c1_31_7),.b(c1_31_6),.c(c1_31_5),.s(s2_32_6),.co(c2_32_6)
);
wire c2_32_7, s2_32_7;
full_adder fa2_32_7 (
.a(c1_31_4),.b(c1_31_3),.c(c1_31_2),.s(s2_32_7),.co(c2_32_7)
);
wire c2_33_1, s2_33_1;
full_adder fa2_33_1 (
.a(s1_33_10),.b(s1_33_9),.c(s1_33_8),.s(s2_33_1),.co(c2_33_1)
);
wire c2_33_2, s2_33_2;
full_adder fa2_33_2 (
.a(s1_33_7),.b(s1_33_6),.c(s1_33_5),.s(s2_33_2),.co(c2_33_2)
);
wire c2_33_3, s2_33_3;
full_adder fa2_33_3 (
.a(s1_33_4),.b(s1_33_3),.c(s1_33_2),.s(s2_33_3),.co(c2_33_3)
);
wire c2_33_4, s2_33_4;
full_adder fa2_33_4 (
.a(s1_33_1),.b(c1_32_10),.c(c1_32_9),.s(s2_33_4),.co(c2_33_4)
);
wire c2_33_5, s2_33_5;
full_adder fa2_33_5 (
.a(c1_32_8),.b(c1_32_7),.c(c1_32_6),.s(s2_33_5),.co(c2_33_5)
);
wire c2_33_6, s2_33_6;
full_adder fa2_33_6 (
.a(c1_32_5),.b(c1_32_4),.c(c1_32_3),.s(s2_33_6),.co(c2_33_6)
);
wire c2_33_7, s2_33_7;
half_adder ha2_33_7 (
.a(c1_32_2),.b(c1_32_1),.p(s2_33_7),.g(c2_33_7)
);
wire c2_34_1, s2_34_1;
full_adder fa2_34_1 (
.a(s1_34_10),.b(s1_34_9),.c(s1_34_8),.s(s2_34_1),.co(c2_34_1)
);
wire c2_34_2, s2_34_2;
full_adder fa2_34_2 (
.a(s1_34_7),.b(s1_34_6),.c(s1_34_5),.s(s2_34_2),.co(c2_34_2)
);
wire c2_34_3, s2_34_3;
full_adder fa2_34_3 (
.a(s1_34_4),.b(s1_34_3),.c(s1_34_2),.s(s2_34_3),.co(c2_34_3)
);
wire c2_34_4, s2_34_4;
full_adder fa2_34_4 (
.a(s1_34_1),.b(c1_33_10),.c(c1_33_9),.s(s2_34_4),.co(c2_34_4)
);
wire c2_34_5, s2_34_5;
full_adder fa2_34_5 (
.a(c1_33_8),.b(c1_33_7),.c(c1_33_6),.s(s2_34_5),.co(c2_34_5)
);
wire c2_34_6, s2_34_6;
full_adder fa2_34_6 (
.a(c1_33_5),.b(c1_33_4),.c(c1_33_3),.s(s2_34_6),.co(c2_34_6)
);
wire c2_34_7, s2_34_7;
half_adder ha2_34_7 (
.a(c1_33_2),.b(c1_33_1),.p(s2_34_7),.g(c2_34_7)
);
wire c2_35_1, s2_35_1;
full_adder fa2_35_1 (
.a(A[31] & B[4]),.b(s1_35_9),.c(s1_35_8),.s(s2_35_1),.co(c2_35_1)
);
wire c2_35_2, s2_35_2;
full_adder fa2_35_2 (
.a(s1_35_7),.b(s1_35_6),.c(s1_35_5),.s(s2_35_2),.co(c2_35_2)
);
wire c2_35_3, s2_35_3;
full_adder fa2_35_3 (
.a(s1_35_4),.b(s1_35_3),.c(s1_35_2),.s(s2_35_3),.co(c2_35_3)
);
wire c2_35_4, s2_35_4;
full_adder fa2_35_4 (
.a(s1_35_1),.b(c1_34_10),.c(c1_34_9),.s(s2_35_4),.co(c2_35_4)
);
wire c2_35_5, s2_35_5;
full_adder fa2_35_5 (
.a(c1_34_8),.b(c1_34_7),.c(c1_34_6),.s(s2_35_5),.co(c2_35_5)
);
wire c2_35_6, s2_35_6;
full_adder fa2_35_6 (
.a(c1_34_5),.b(c1_34_4),.c(c1_34_3),.s(s2_35_6),.co(c2_35_6)
);
wire c2_35_7, s2_35_7;
half_adder ha2_35_7 (
.a(c1_34_2),.b(c1_34_1),.p(s2_35_7),.g(c2_35_7)
);
wire c2_36_1, s2_36_1;
full_adder fa2_36_1 (
.a(s1_36_9),.b(s1_36_8),.c(s1_36_7),.s(s2_36_1),.co(c2_36_1)
);
wire c2_36_2, s2_36_2;
full_adder fa2_36_2 (
.a(s1_36_6),.b(s1_36_5),.c(s1_36_4),.s(s2_36_2),.co(c2_36_2)
);
wire c2_36_3, s2_36_3;
full_adder fa2_36_3 (
.a(s1_36_3),.b(s1_36_2),.c(s1_36_1),.s(s2_36_3),.co(c2_36_3)
);
wire c2_36_4, s2_36_4;
full_adder fa2_36_4 (
.a(c1_35_9),.b(c1_35_8),.c(c1_35_7),.s(s2_36_4),.co(c2_36_4)
);
wire c2_36_5, s2_36_5;
full_adder fa2_36_5 (
.a(c1_35_6),.b(c1_35_5),.c(c1_35_4),.s(s2_36_5),.co(c2_36_5)
);
wire c2_36_6, s2_36_6;
full_adder fa2_36_6 (
.a(c1_35_3),.b(c1_35_2),.c(c1_35_1),.s(s2_36_6),.co(c2_36_6)
);
wire c2_37_1, s2_37_1;
full_adder fa2_37_1 (
.a(s1_37_9),.b(s1_37_8),.c(s1_37_7),.s(s2_37_1),.co(c2_37_1)
);
wire c2_37_2, s2_37_2;
full_adder fa2_37_2 (
.a(s1_37_6),.b(s1_37_5),.c(s1_37_4),.s(s2_37_2),.co(c2_37_2)
);
wire c2_37_3, s2_37_3;
full_adder fa2_37_3 (
.a(s1_37_3),.b(s1_37_2),.c(s1_37_1),.s(s2_37_3),.co(c2_37_3)
);
wire c2_37_4, s2_37_4;
full_adder fa2_37_4 (
.a(c1_36_9),.b(c1_36_8),.c(c1_36_7),.s(s2_37_4),.co(c2_37_4)
);
wire c2_37_5, s2_37_5;
full_adder fa2_37_5 (
.a(c1_36_6),.b(c1_36_5),.c(c1_36_4),.s(s2_37_5),.co(c2_37_5)
);
wire c2_37_6, s2_37_6;
full_adder fa2_37_6 (
.a(c1_36_3),.b(c1_36_2),.c(c1_36_1),.s(s2_37_6),.co(c2_37_6)
);
wire c2_38_1, s2_38_1;
full_adder fa2_38_1 (
.a(A[31] & B[7]),.b(s1_38_8),.c(s1_38_7),.s(s2_38_1),.co(c2_38_1)
);
wire c2_38_2, s2_38_2;
full_adder fa2_38_2 (
.a(s1_38_6),.b(s1_38_5),.c(s1_38_4),.s(s2_38_2),.co(c2_38_2)
);
wire c2_38_3, s2_38_3;
full_adder fa2_38_3 (
.a(s1_38_3),.b(s1_38_2),.c(s1_38_1),.s(s2_38_3),.co(c2_38_3)
);
wire c2_38_4, s2_38_4;
full_adder fa2_38_4 (
.a(c1_37_9),.b(c1_37_8),.c(c1_37_7),.s(s2_38_4),.co(c2_38_4)
);
wire c2_38_5, s2_38_5;
full_adder fa2_38_5 (
.a(c1_37_6),.b(c1_37_5),.c(c1_37_4),.s(s2_38_5),.co(c2_38_5)
);
wire c2_38_6, s2_38_6;
full_adder fa2_38_6 (
.a(c1_37_3),.b(c1_37_2),.c(c1_37_1),.s(s2_38_6),.co(c2_38_6)
);
wire c2_39_1, s2_39_1;
full_adder fa2_39_1 (
.a(s1_39_8),.b(s1_39_7),.c(s1_39_6),.s(s2_39_1),.co(c2_39_1)
);
wire c2_39_2, s2_39_2;
full_adder fa2_39_2 (
.a(s1_39_5),.b(s1_39_4),.c(s1_39_3),.s(s2_39_2),.co(c2_39_2)
);
wire c2_39_3, s2_39_3;
full_adder fa2_39_3 (
.a(s1_39_2),.b(s1_39_1),.c(c1_38_8),.s(s2_39_3),.co(c2_39_3)
);
wire c2_39_4, s2_39_4;
full_adder fa2_39_4 (
.a(c1_38_7),.b(c1_38_6),.c(c1_38_5),.s(s2_39_4),.co(c2_39_4)
);
wire c2_39_5, s2_39_5;
full_adder fa2_39_5 (
.a(c1_38_4),.b(c1_38_3),.c(c1_38_2),.s(s2_39_5),.co(c2_39_5)
);
wire c2_40_1, s2_40_1;
full_adder fa2_40_1 (
.a(s1_40_8),.b(s1_40_7),.c(s1_40_6),.s(s2_40_1),.co(c2_40_1)
);
wire c2_40_2, s2_40_2;
full_adder fa2_40_2 (
.a(s1_40_5),.b(s1_40_4),.c(s1_40_3),.s(s2_40_2),.co(c2_40_2)
);
wire c2_40_3, s2_40_3;
full_adder fa2_40_3 (
.a(s1_40_2),.b(s1_40_1),.c(c1_39_8),.s(s2_40_3),.co(c2_40_3)
);
wire c2_40_4, s2_40_4;
full_adder fa2_40_4 (
.a(c1_39_7),.b(c1_39_6),.c(c1_39_5),.s(s2_40_4),.co(c2_40_4)
);
wire c2_40_5, s2_40_5;
full_adder fa2_40_5 (
.a(c1_39_4),.b(c1_39_3),.c(c1_39_2),.s(s2_40_5),.co(c2_40_5)
);
wire c2_41_1, s2_41_1;
full_adder fa2_41_1 (
.a(A[31] & B[10]),.b(s1_41_7),.c(s1_41_6),.s(s2_41_1),.co(c2_41_1)
);
wire c2_41_2, s2_41_2;
full_adder fa2_41_2 (
.a(s1_41_5),.b(s1_41_4),.c(s1_41_3),.s(s2_41_2),.co(c2_41_2)
);
wire c2_41_3, s2_41_3;
full_adder fa2_41_3 (
.a(s1_41_2),.b(s1_41_1),.c(c1_40_8),.s(s2_41_3),.co(c2_41_3)
);
wire c2_41_4, s2_41_4;
full_adder fa2_41_4 (
.a(c1_40_7),.b(c1_40_6),.c(c1_40_5),.s(s2_41_4),.co(c2_41_4)
);
wire c2_41_5, s2_41_5;
full_adder fa2_41_5 (
.a(c1_40_4),.b(c1_40_3),.c(c1_40_2),.s(s2_41_5),.co(c2_41_5)
);
wire c2_42_1, s2_42_1;
full_adder fa2_42_1 (
.a(s1_42_7),.b(s1_42_6),.c(s1_42_5),.s(s2_42_1),.co(c2_42_1)
);
wire c2_42_2, s2_42_2;
full_adder fa2_42_2 (
.a(s1_42_4),.b(s1_42_3),.c(s1_42_2),.s(s2_42_2),.co(c2_42_2)
);
wire c2_42_3, s2_42_3;
full_adder fa2_42_3 (
.a(s1_42_1),.b(c1_41_7),.c(c1_41_6),.s(s2_42_3),.co(c2_42_3)
);
wire c2_42_4, s2_42_4;
full_adder fa2_42_4 (
.a(c1_41_5),.b(c1_41_4),.c(c1_41_3),.s(s2_42_4),.co(c2_42_4)
);
wire c2_42_5, s2_42_5;
half_adder ha2_42_5 (
.a(c1_41_2),.b(c1_41_1),.p(s2_42_5),.g(c2_42_5)
);
wire c2_43_1, s2_43_1;
full_adder fa2_43_1 (
.a(s1_43_7),.b(s1_43_6),.c(s1_43_5),.s(s2_43_1),.co(c2_43_1)
);
wire c2_43_2, s2_43_2;
full_adder fa2_43_2 (
.a(s1_43_4),.b(s1_43_3),.c(s1_43_2),.s(s2_43_2),.co(c2_43_2)
);
wire c2_43_3, s2_43_3;
full_adder fa2_43_3 (
.a(s1_43_1),.b(c1_42_7),.c(c1_42_6),.s(s2_43_3),.co(c2_43_3)
);
wire c2_43_4, s2_43_4;
full_adder fa2_43_4 (
.a(c1_42_5),.b(c1_42_4),.c(c1_42_3),.s(s2_43_4),.co(c2_43_4)
);
wire c2_43_5, s2_43_5;
half_adder ha2_43_5 (
.a(c1_42_2),.b(c1_42_1),.p(s2_43_5),.g(c2_43_5)
);
wire c2_44_1, s2_44_1;
full_adder fa2_44_1 (
.a(A[31] & B[13]),.b(s1_44_6),.c(s1_44_5),.s(s2_44_1),.co(c2_44_1)
);
wire c2_44_2, s2_44_2;
full_adder fa2_44_2 (
.a(s1_44_4),.b(s1_44_3),.c(s1_44_2),.s(s2_44_2),.co(c2_44_2)
);
wire c2_44_3, s2_44_3;
full_adder fa2_44_3 (
.a(s1_44_1),.b(c1_43_7),.c(c1_43_6),.s(s2_44_3),.co(c2_44_3)
);
wire c2_44_4, s2_44_4;
full_adder fa2_44_4 (
.a(c1_43_5),.b(c1_43_4),.c(c1_43_3),.s(s2_44_4),.co(c2_44_4)
);
wire c2_44_5, s2_44_5;
half_adder ha2_44_5 (
.a(c1_43_2),.b(c1_43_1),.p(s2_44_5),.g(c2_44_5)
);
wire c2_45_1, s2_45_1;
full_adder fa2_45_1 (
.a(s1_45_6),.b(s1_45_5),.c(s1_45_4),.s(s2_45_1),.co(c2_45_1)
);
wire c2_45_2, s2_45_2;
full_adder fa2_45_2 (
.a(s1_45_3),.b(s1_45_2),.c(s1_45_1),.s(s2_45_2),.co(c2_45_2)
);
wire c2_45_3, s2_45_3;
full_adder fa2_45_3 (
.a(c1_44_6),.b(c1_44_5),.c(c1_44_4),.s(s2_45_3),.co(c2_45_3)
);
wire c2_45_4, s2_45_4;
full_adder fa2_45_4 (
.a(c1_44_3),.b(c1_44_2),.c(c1_44_1),.s(s2_45_4),.co(c2_45_4)
);
wire c2_46_1, s2_46_1;
full_adder fa2_46_1 (
.a(s1_46_6),.b(s1_46_5),.c(s1_46_4),.s(s2_46_1),.co(c2_46_1)
);
wire c2_46_2, s2_46_2;
full_adder fa2_46_2 (
.a(s1_46_3),.b(s1_46_2),.c(s1_46_1),.s(s2_46_2),.co(c2_46_2)
);
wire c2_46_3, s2_46_3;
full_adder fa2_46_3 (
.a(c1_45_6),.b(c1_45_5),.c(c1_45_4),.s(s2_46_3),.co(c2_46_3)
);
wire c2_46_4, s2_46_4;
full_adder fa2_46_4 (
.a(c1_45_3),.b(c1_45_2),.c(c1_45_1),.s(s2_46_4),.co(c2_46_4)
);
wire c2_47_1, s2_47_1;
full_adder fa2_47_1 (
.a(A[31] & B[16]),.b(s1_47_5),.c(s1_47_4),.s(s2_47_1),.co(c2_47_1)
);
wire c2_47_2, s2_47_2;
full_adder fa2_47_2 (
.a(s1_47_3),.b(s1_47_2),.c(s1_47_1),.s(s2_47_2),.co(c2_47_2)
);
wire c2_47_3, s2_47_3;
full_adder fa2_47_3 (
.a(c1_46_6),.b(c1_46_5),.c(c1_46_4),.s(s2_47_3),.co(c2_47_3)
);
wire c2_47_4, s2_47_4;
full_adder fa2_47_4 (
.a(c1_46_3),.b(c1_46_2),.c(c1_46_1),.s(s2_47_4),.co(c2_47_4)
);
wire c2_48_1, s2_48_1;
full_adder fa2_48_1 (
.a(s1_48_5),.b(s1_48_4),.c(s1_48_3),.s(s2_48_1),.co(c2_48_1)
);
wire c2_48_2, s2_48_2;
full_adder fa2_48_2 (
.a(s1_48_2),.b(s1_48_1),.c(c1_47_5),.s(s2_48_2),.co(c2_48_2)
);
wire c2_48_3, s2_48_3;
full_adder fa2_48_3 (
.a(c1_47_4),.b(c1_47_3),.c(c1_47_2),.s(s2_48_3),.co(c2_48_3)
);
wire c2_49_1, s2_49_1;
full_adder fa2_49_1 (
.a(s1_49_5),.b(s1_49_4),.c(s1_49_3),.s(s2_49_1),.co(c2_49_1)
);
wire c2_49_2, s2_49_2;
full_adder fa2_49_2 (
.a(s1_49_2),.b(s1_49_1),.c(c1_48_5),.s(s2_49_2),.co(c2_49_2)
);
wire c2_49_3, s2_49_3;
full_adder fa2_49_3 (
.a(c1_48_4),.b(c1_48_3),.c(c1_48_2),.s(s2_49_3),.co(c2_49_3)
);
wire c2_50_1, s2_50_1;
full_adder fa2_50_1 (
.a(A[31] & B[19]),.b(s1_50_4),.c(s1_50_3),.s(s2_50_1),.co(c2_50_1)
);
wire c2_50_2, s2_50_2;
full_adder fa2_50_2 (
.a(s1_50_2),.b(s1_50_1),.c(c1_49_5),.s(s2_50_2),.co(c2_50_2)
);
wire c2_50_3, s2_50_3;
full_adder fa2_50_3 (
.a(c1_49_4),.b(c1_49_3),.c(c1_49_2),.s(s2_50_3),.co(c2_50_3)
);
wire c2_51_1, s2_51_1;
full_adder fa2_51_1 (
.a(s1_51_4),.b(s1_51_3),.c(s1_51_2),.s(s2_51_1),.co(c2_51_1)
);
wire c2_51_2, s2_51_2;
full_adder fa2_51_2 (
.a(s1_51_1),.b(c1_50_4),.c(c1_50_3),.s(s2_51_2),.co(c2_51_2)
);
wire c2_51_3, s2_51_3;
half_adder ha2_51_3 (
.a(c1_50_2),.b(c1_50_1),.p(s2_51_3),.g(c2_51_3)
);
wire c2_52_1, s2_52_1;
full_adder fa2_52_1 (
.a(s1_52_4),.b(s1_52_3),.c(s1_52_2),.s(s2_52_1),.co(c2_52_1)
);
wire c2_52_2, s2_52_2;
full_adder fa2_52_2 (
.a(s1_52_1),.b(c1_51_4),.c(c1_51_3),.s(s2_52_2),.co(c2_52_2)
);
wire c2_52_3, s2_52_3;
half_adder ha2_52_3 (
.a(c1_51_2),.b(c1_51_1),.p(s2_52_3),.g(c2_52_3)
);
wire c2_53_1, s2_53_1;
full_adder fa2_53_1 (
.a(A[31] & B[22]),.b(s1_53_3),.c(s1_53_2),.s(s2_53_1),.co(c2_53_1)
);
wire c2_53_2, s2_53_2;
full_adder fa2_53_2 (
.a(s1_53_1),.b(c1_52_4),.c(c1_52_3),.s(s2_53_2),.co(c2_53_2)
);
wire c2_53_3, s2_53_3;
half_adder ha2_53_3 (
.a(c1_52_2),.b(c1_52_1),.p(s2_53_3),.g(c2_53_3)
);
wire c2_54_1, s2_54_1;
full_adder fa2_54_1 (
.a(s1_54_3),.b(s1_54_2),.c(s1_54_1),.s(s2_54_1),.co(c2_54_1)
);
wire c2_54_2, s2_54_2;
full_adder fa2_54_2 (
.a(c1_53_3),.b(c1_53_2),.c(c1_53_1),.s(s2_54_2),.co(c2_54_2)
);
wire c2_55_1, s2_55_1;
full_adder fa2_55_1 (
.a(s1_55_3),.b(s1_55_2),.c(s1_55_1),.s(s2_55_1),.co(c2_55_1)
);
wire c2_55_2, s2_55_2;
full_adder fa2_55_2 (
.a(c1_54_3),.b(c1_54_2),.c(c1_54_1),.s(s2_55_2),.co(c2_55_2)
);
wire c2_56_1, s2_56_1;
full_adder fa2_56_1 (
.a(A[31] & B[25]),.b(s1_56_2),.c(s1_56_1),.s(s2_56_1),.co(c2_56_1)
);
wire c2_56_2, s2_56_2;
full_adder fa2_56_2 (
.a(c1_55_3),.b(c1_55_2),.c(c1_55_1),.s(s2_56_2),.co(c2_56_2)
);
wire c2_57_1, s2_57_1;
full_adder fa2_57_1 (
.a(s1_57_2),.b(s1_57_1),.c(c1_56_2),.s(s2_57_1),.co(c2_57_1)
);
wire c2_58_1, s2_58_1;
full_adder fa2_58_1 (
.a(s1_58_2),.b(s1_58_1),.c(c1_57_2),.s(s2_58_1),.co(c2_58_1)
);
wire c2_59_1, s2_59_1;
full_adder fa2_59_1 (
.a(A[31] & B[28]),.b(s1_59_1),.c(c1_58_2),.s(s2_59_1),.co(c2_59_1)
);
wire c2_60_1, s2_60_1;
half_adder ha2_60_1 (
.a(s1_60_1),.b(c1_59_1),.p(s2_60_1),.g(c2_60_1)
);
wire c2_61_1, s2_61_1;
half_adder ha2_61_1 (
.a(s1_61_1),.b(c1_60_1),.p(s2_61_1),.g(c2_61_1)
);
wire c2_62_1, s2_62_1;
half_adder ha2_62_1 (
.a(A[31] & B[31]),.b(c1_61_1),.p(s2_62_1),.g(c2_62_1)
);
wire c3_3_1, s3_3_1;
half_adder ha3_3_1 (
.a(s2_3_1),.b(c2_2_1),.p(s3_3_1),.g(c3_3_1)
);
wire c3_4_1, s3_4_1;
half_adder ha3_4_1 (
.a(s2_4_1),.b(c2_3_1),.p(s3_4_1),.g(c3_4_1)
);
wire c3_5_1, s3_5_1;
full_adder fa3_5_1 (
.a(c1_4_1),.b(s2_5_1),.c(c2_4_1),.s(s3_5_1),.co(c3_5_1)
);
wire c3_6_1, s3_6_1;
full_adder fa3_6_1 (
.a(s2_6_2),.b(s2_6_1),.c(c2_5_1),.s(s3_6_1),.co(c3_6_1)
);
wire c3_7_1, s3_7_1;
full_adder fa3_7_1 (
.a(s2_7_2),.b(s2_7_1),.c(c2_6_2),.s(s3_7_1),.co(c3_7_1)
);
wire c3_8_1, s3_8_1;
full_adder fa3_8_1 (
.a(s2_8_2),.b(s2_8_1),.c(c2_7_2),.s(s3_8_1),.co(c3_8_1)
);
wire c3_9_1, s3_9_1;
full_adder fa3_9_1 (
.a(c1_8_1),.b(s2_9_2),.c(s2_9_1),.s(s3_9_1),.co(c3_9_1)
);
wire c3_9_2, s3_9_2;
half_adder ha3_9_2 (
.a(c2_8_2),.b(c2_8_1),.p(s3_9_2),.g(c3_9_2)
);
wire c3_10_1, s3_10_1;
full_adder fa3_10_1 (
.a(c1_9_1),.b(s2_10_2),.c(s2_10_1),.s(s3_10_1),.co(c3_10_1)
);
wire c3_10_2, s3_10_2;
half_adder ha3_10_2 (
.a(c2_9_2),.b(c2_9_1),.p(s3_10_2),.g(c3_10_2)
);
wire c3_11_1, s3_11_1;
full_adder fa3_11_1 (
.a(s2_11_3),.b(s2_11_2),.c(s2_11_1),.s(s3_11_1),.co(c3_11_1)
);
wire c3_11_2, s3_11_2;
half_adder ha3_11_2 (
.a(c2_10_2),.b(c2_10_1),.p(s3_11_2),.g(c3_11_2)
);
wire c3_12_1, s3_12_1;
full_adder fa3_12_1 (
.a(s2_12_3),.b(s2_12_2),.c(s2_12_1),.s(s3_12_1),.co(c3_12_1)
);
wire c3_12_2, s3_12_2;
full_adder fa3_12_2 (
.a(c2_11_3),.b(c2_11_2),.c(c2_11_1),.s(s3_12_2),.co(c3_12_2)
);
wire c3_13_1, s3_13_1;
full_adder fa3_13_1 (
.a(s2_13_3),.b(s2_13_2),.c(s2_13_1),.s(s3_13_1),.co(c3_13_1)
);
wire c3_13_2, s3_13_2;
full_adder fa3_13_2 (
.a(c2_12_3),.b(c2_12_2),.c(c2_12_1),.s(s3_13_2),.co(c3_13_2)
);
wire c3_14_1, s3_14_1;
full_adder fa3_14_1 (
.a(c1_13_1),.b(s2_14_3),.c(s2_14_2),.s(s3_14_1),.co(c3_14_1)
);
wire c3_14_2, s3_14_2;
full_adder fa3_14_2 (
.a(s2_14_1),.b(c2_13_3),.c(c2_13_2),.s(s3_14_2),.co(c3_14_2)
);
wire c3_15_1, s3_15_1;
full_adder fa3_15_1 (
.a(s2_15_4),.b(s2_15_3),.c(s2_15_2),.s(s3_15_1),.co(c3_15_1)
);
wire c3_15_2, s3_15_2;
full_adder fa3_15_2 (
.a(s2_15_1),.b(c2_14_3),.c(c2_14_2),.s(s3_15_2),.co(c3_15_2)
);
wire c3_16_1, s3_16_1;
full_adder fa3_16_1 (
.a(s2_16_4),.b(s2_16_3),.c(s2_16_2),.s(s3_16_1),.co(c3_16_1)
);
wire c3_16_2, s3_16_2;
full_adder fa3_16_2 (
.a(s2_16_1),.b(c2_15_4),.c(c2_15_3),.s(s3_16_2),.co(c3_16_2)
);
wire c3_16_3, s3_16_3;
half_adder ha3_16_3 (
.a(c2_15_2),.b(c2_15_1),.p(s3_16_3),.g(c3_16_3)
);
wire c3_17_1, s3_17_1;
full_adder fa3_17_1 (
.a(s2_17_4),.b(s2_17_3),.c(s2_17_2),.s(s3_17_1),.co(c3_17_1)
);
wire c3_17_2, s3_17_2;
full_adder fa3_17_2 (
.a(s2_17_1),.b(c2_16_4),.c(c2_16_3),.s(s3_17_2),.co(c3_17_2)
);
wire c3_17_3, s3_17_3;
half_adder ha3_17_3 (
.a(c2_16_2),.b(c2_16_1),.p(s3_17_3),.g(c3_17_3)
);
wire c3_18_1, s3_18_1;
full_adder fa3_18_1 (
.a(c1_17_1),.b(s2_18_4),.c(s2_18_3),.s(s3_18_1),.co(c3_18_1)
);
wire c3_18_2, s3_18_2;
full_adder fa3_18_2 (
.a(s2_18_2),.b(s2_18_1),.c(c2_17_4),.s(s3_18_2),.co(c3_18_2)
);
wire c3_18_3, s3_18_3;
full_adder fa3_18_3 (
.a(c2_17_3),.b(c2_17_2),.c(c2_17_1),.s(s3_18_3),.co(c3_18_3)
);
wire c3_19_1, s3_19_1;
full_adder fa3_19_1 (
.a(c1_18_1),.b(s2_19_4),.c(s2_19_3),.s(s3_19_1),.co(c3_19_1)
);
wire c3_19_2, s3_19_2;
full_adder fa3_19_2 (
.a(s2_19_2),.b(s2_19_1),.c(c2_18_4),.s(s3_19_2),.co(c3_19_2)
);
wire c3_19_3, s3_19_3;
full_adder fa3_19_3 (
.a(c2_18_3),.b(c2_18_2),.c(c2_18_1),.s(s3_19_3),.co(c3_19_3)
);
wire c3_20_1, s3_20_1;
full_adder fa3_20_1 (
.a(s2_20_5),.b(s2_20_4),.c(s2_20_3),.s(s3_20_1),.co(c3_20_1)
);
wire c3_20_2, s3_20_2;
full_adder fa3_20_2 (
.a(s2_20_2),.b(s2_20_1),.c(c2_19_4),.s(s3_20_2),.co(c3_20_2)
);
wire c3_20_3, s3_20_3;
full_adder fa3_20_3 (
.a(c2_19_3),.b(c2_19_2),.c(c2_19_1),.s(s3_20_3),.co(c3_20_3)
);
wire c3_21_1, s3_21_1;
full_adder fa3_21_1 (
.a(s2_21_5),.b(s2_21_4),.c(s2_21_3),.s(s3_21_1),.co(c3_21_1)
);
wire c3_21_2, s3_21_2;
full_adder fa3_21_2 (
.a(s2_21_2),.b(s2_21_1),.c(c2_20_5),.s(s3_21_2),.co(c3_21_2)
);
wire c3_21_3, s3_21_3;
full_adder fa3_21_3 (
.a(c2_20_4),.b(c2_20_3),.c(c2_20_2),.s(s3_21_3),.co(c3_21_3)
);
wire c3_22_1, s3_22_1;
full_adder fa3_22_1 (
.a(s2_22_5),.b(s2_22_4),.c(s2_22_3),.s(s3_22_1),.co(c3_22_1)
);
wire c3_22_2, s3_22_2;
full_adder fa3_22_2 (
.a(s2_22_2),.b(s2_22_1),.c(c2_21_5),.s(s3_22_2),.co(c3_22_2)
);
wire c3_22_3, s3_22_3;
full_adder fa3_22_3 (
.a(c2_21_4),.b(c2_21_3),.c(c2_21_2),.s(s3_22_3),.co(c3_22_3)
);
wire c3_23_1, s3_23_1;
full_adder fa3_23_1 (
.a(c1_22_1),.b(s2_23_5),.c(s2_23_4),.s(s3_23_1),.co(c3_23_1)
);
wire c3_23_2, s3_23_2;
full_adder fa3_23_2 (
.a(s2_23_3),.b(s2_23_2),.c(s2_23_1),.s(s3_23_2),.co(c3_23_2)
);
wire c3_23_3, s3_23_3;
full_adder fa3_23_3 (
.a(c2_22_5),.b(c2_22_4),.c(c2_22_3),.s(s3_23_3),.co(c3_23_3)
);
wire c3_23_4, s3_23_4;
half_adder ha3_23_4 (
.a(c2_22_2),.b(c2_22_1),.p(s3_23_4),.g(c3_23_4)
);
wire c3_24_1, s3_24_1;
full_adder fa3_24_1 (
.a(s2_24_6),.b(s2_24_5),.c(s2_24_4),.s(s3_24_1),.co(c3_24_1)
);
wire c3_24_2, s3_24_2;
full_adder fa3_24_2 (
.a(s2_24_3),.b(s2_24_2),.c(s2_24_1),.s(s3_24_2),.co(c3_24_2)
);
wire c3_24_3, s3_24_3;
full_adder fa3_24_3 (
.a(c2_23_5),.b(c2_23_4),.c(c2_23_3),.s(s3_24_3),.co(c3_24_3)
);
wire c3_24_4, s3_24_4;
half_adder ha3_24_4 (
.a(c2_23_2),.b(c2_23_1),.p(s3_24_4),.g(c3_24_4)
);
wire c3_25_1, s3_25_1;
full_adder fa3_25_1 (
.a(s2_25_6),.b(s2_25_5),.c(s2_25_4),.s(s3_25_1),.co(c3_25_1)
);
wire c3_25_2, s3_25_2;
full_adder fa3_25_2 (
.a(s2_25_3),.b(s2_25_2),.c(s2_25_1),.s(s3_25_2),.co(c3_25_2)
);
wire c3_25_3, s3_25_3;
full_adder fa3_25_3 (
.a(c2_24_6),.b(c2_24_5),.c(c2_24_4),.s(s3_25_3),.co(c3_25_3)
);
wire c3_25_4, s3_25_4;
full_adder fa3_25_4 (
.a(c2_24_3),.b(c2_24_2),.c(c2_24_1),.s(s3_25_4),.co(c3_25_4)
);
wire c3_26_1, s3_26_1;
full_adder fa3_26_1 (
.a(s2_26_6),.b(s2_26_5),.c(s2_26_4),.s(s3_26_1),.co(c3_26_1)
);
wire c3_26_2, s3_26_2;
full_adder fa3_26_2 (
.a(s2_26_3),.b(s2_26_2),.c(s2_26_1),.s(s3_26_2),.co(c3_26_2)
);
wire c3_26_3, s3_26_3;
full_adder fa3_26_3 (
.a(c2_25_6),.b(c2_25_5),.c(c2_25_4),.s(s3_26_3),.co(c3_26_3)
);
wire c3_26_4, s3_26_4;
full_adder fa3_26_4 (
.a(c2_25_3),.b(c2_25_2),.c(c2_25_1),.s(s3_26_4),.co(c3_26_4)
);
wire c3_27_1, s3_27_1;
full_adder fa3_27_1 (
.a(c1_26_1),.b(s2_27_6),.c(s2_27_5),.s(s3_27_1),.co(c3_27_1)
);
wire c3_27_2, s3_27_2;
full_adder fa3_27_2 (
.a(s2_27_4),.b(s2_27_3),.c(s2_27_2),.s(s3_27_2),.co(c3_27_2)
);
wire c3_27_3, s3_27_3;
full_adder fa3_27_3 (
.a(s2_27_1),.b(c2_26_6),.c(c2_26_5),.s(s3_27_3),.co(c3_27_3)
);
wire c3_27_4, s3_27_4;
full_adder fa3_27_4 (
.a(c2_26_4),.b(c2_26_3),.c(c2_26_2),.s(s3_27_4),.co(c3_27_4)
);
wire c3_28_1, s3_28_1;
full_adder fa3_28_1 (
.a(c1_27_1),.b(s2_28_6),.c(s2_28_5),.s(s3_28_1),.co(c3_28_1)
);
wire c3_28_2, s3_28_2;
full_adder fa3_28_2 (
.a(s2_28_4),.b(s2_28_3),.c(s2_28_2),.s(s3_28_2),.co(c3_28_2)
);
wire c3_28_3, s3_28_3;
full_adder fa3_28_3 (
.a(s2_28_1),.b(c2_27_6),.c(c2_27_5),.s(s3_28_3),.co(c3_28_3)
);
wire c3_28_4, s3_28_4;
full_adder fa3_28_4 (
.a(c2_27_4),.b(c2_27_3),.c(c2_27_2),.s(s3_28_4),.co(c3_28_4)
);
wire c3_29_1, s3_29_1;
full_adder fa3_29_1 (
.a(s2_29_7),.b(s2_29_6),.c(s2_29_5),.s(s3_29_1),.co(c3_29_1)
);
wire c3_29_2, s3_29_2;
full_adder fa3_29_2 (
.a(s2_29_4),.b(s2_29_3),.c(s2_29_2),.s(s3_29_2),.co(c3_29_2)
);
wire c3_29_3, s3_29_3;
full_adder fa3_29_3 (
.a(s2_29_1),.b(c2_28_6),.c(c2_28_5),.s(s3_29_3),.co(c3_29_3)
);
wire c3_29_4, s3_29_4;
full_adder fa3_29_4 (
.a(c2_28_4),.b(c2_28_3),.c(c2_28_2),.s(s3_29_4),.co(c3_29_4)
);
wire c3_30_1, s3_30_1;
full_adder fa3_30_1 (
.a(s2_30_7),.b(s2_30_6),.c(s2_30_5),.s(s3_30_1),.co(c3_30_1)
);
wire c3_30_2, s3_30_2;
full_adder fa3_30_2 (
.a(s2_30_4),.b(s2_30_3),.c(s2_30_2),.s(s3_30_2),.co(c3_30_2)
);
wire c3_30_3, s3_30_3;
full_adder fa3_30_3 (
.a(s2_30_1),.b(c2_29_7),.c(c2_29_6),.s(s3_30_3),.co(c3_30_3)
);
wire c3_30_4, s3_30_4;
full_adder fa3_30_4 (
.a(c2_29_5),.b(c2_29_4),.c(c2_29_3),.s(s3_30_4),.co(c3_30_4)
);
wire c3_30_5, s3_30_5;
half_adder ha3_30_5 (
.a(c2_29_2),.b(c2_29_1),.p(s3_30_5),.g(c3_30_5)
);
wire c3_31_1, s3_31_1;
full_adder fa3_31_1 (
.a(s2_31_7),.b(s2_31_6),.c(s2_31_5),.s(s3_31_1),.co(c3_31_1)
);
wire c3_31_2, s3_31_2;
full_adder fa3_31_2 (
.a(s2_31_4),.b(s2_31_3),.c(s2_31_2),.s(s3_31_2),.co(c3_31_2)
);
wire c3_31_3, s3_31_3;
full_adder fa3_31_3 (
.a(s2_31_1),.b(c2_30_7),.c(c2_30_6),.s(s3_31_3),.co(c3_31_3)
);
wire c3_31_4, s3_31_4;
full_adder fa3_31_4 (
.a(c2_30_5),.b(c2_30_4),.c(c2_30_3),.s(s3_31_4),.co(c3_31_4)
);
wire c3_31_5, s3_31_5;
half_adder ha3_31_5 (
.a(c2_30_2),.b(c2_30_1),.p(s3_31_5),.g(c3_31_5)
);
wire c3_32_1, s3_32_1;
full_adder fa3_32_1 (
.a(c1_31_1),.b(s2_32_7),.c(s2_32_6),.s(s3_32_1),.co(c3_32_1)
);
wire c3_32_2, s3_32_2;
full_adder fa3_32_2 (
.a(s2_32_5),.b(s2_32_4),.c(s2_32_3),.s(s3_32_2),.co(c3_32_2)
);
wire c3_32_3, s3_32_3;
full_adder fa3_32_3 (
.a(s2_32_2),.b(s2_32_1),.c(c2_31_7),.s(s3_32_3),.co(c3_32_3)
);
wire c3_32_4, s3_32_4;
full_adder fa3_32_4 (
.a(c2_31_6),.b(c2_31_5),.c(c2_31_4),.s(s3_32_4),.co(c3_32_4)
);
wire c3_32_5, s3_32_5;
full_adder fa3_32_5 (
.a(c2_31_3),.b(c2_31_2),.c(c2_31_1),.s(s3_32_5),.co(c3_32_5)
);
wire c3_33_1, s3_33_1;
full_adder fa3_33_1 (
.a(s2_33_7),.b(s2_33_6),.c(s2_33_5),.s(s3_33_1),.co(c3_33_1)
);
wire c3_33_2, s3_33_2;
full_adder fa3_33_2 (
.a(s2_33_4),.b(s2_33_3),.c(s2_33_2),.s(s3_33_2),.co(c3_33_2)
);
wire c3_33_3, s3_33_3;
full_adder fa3_33_3 (
.a(s2_33_1),.b(c2_32_7),.c(c2_32_6),.s(s3_33_3),.co(c3_33_3)
);
wire c3_33_4, s3_33_4;
full_adder fa3_33_4 (
.a(c2_32_5),.b(c2_32_4),.c(c2_32_3),.s(s3_33_4),.co(c3_33_4)
);
wire c3_33_5, s3_33_5;
half_adder ha3_33_5 (
.a(c2_32_2),.b(c2_32_1),.p(s3_33_5),.g(c3_33_5)
);
wire c3_34_1, s3_34_1;
full_adder fa3_34_1 (
.a(s2_34_7),.b(s2_34_6),.c(s2_34_5),.s(s3_34_1),.co(c3_34_1)
);
wire c3_34_2, s3_34_2;
full_adder fa3_34_2 (
.a(s2_34_4),.b(s2_34_3),.c(s2_34_2),.s(s3_34_2),.co(c3_34_2)
);
wire c3_34_3, s3_34_3;
full_adder fa3_34_3 (
.a(s2_34_1),.b(c2_33_7),.c(c2_33_6),.s(s3_34_3),.co(c3_34_3)
);
wire c3_34_4, s3_34_4;
full_adder fa3_34_4 (
.a(c2_33_5),.b(c2_33_4),.c(c2_33_3),.s(s3_34_4),.co(c3_34_4)
);
wire c3_34_5, s3_34_5;
half_adder ha3_34_5 (
.a(c2_33_2),.b(c2_33_1),.p(s3_34_5),.g(c3_34_5)
);
wire c3_35_1, s3_35_1;
full_adder fa3_35_1 (
.a(s2_35_7),.b(s2_35_6),.c(s2_35_5),.s(s3_35_1),.co(c3_35_1)
);
wire c3_35_2, s3_35_2;
full_adder fa3_35_2 (
.a(s2_35_4),.b(s2_35_3),.c(s2_35_2),.s(s3_35_2),.co(c3_35_2)
);
wire c3_35_3, s3_35_3;
full_adder fa3_35_3 (
.a(s2_35_1),.b(c2_34_7),.c(c2_34_6),.s(s3_35_3),.co(c3_35_3)
);
wire c3_35_4, s3_35_4;
full_adder fa3_35_4 (
.a(c2_34_5),.b(c2_34_4),.c(c2_34_3),.s(s3_35_4),.co(c3_35_4)
);
wire c3_35_5, s3_35_5;
half_adder ha3_35_5 (
.a(c2_34_2),.b(c2_34_1),.p(s3_35_5),.g(c3_35_5)
);
wire c3_36_1, s3_36_1;
full_adder fa3_36_1 (
.a(s2_36_6),.b(s2_36_5),.c(s2_36_4),.s(s3_36_1),.co(c3_36_1)
);
wire c3_36_2, s3_36_2;
full_adder fa3_36_2 (
.a(s2_36_3),.b(s2_36_2),.c(s2_36_1),.s(s3_36_2),.co(c3_36_2)
);
wire c3_36_3, s3_36_3;
full_adder fa3_36_3 (
.a(c2_35_7),.b(c2_35_6),.c(c2_35_5),.s(s3_36_3),.co(c3_36_3)
);
wire c3_36_4, s3_36_4;
full_adder fa3_36_4 (
.a(c2_35_4),.b(c2_35_3),.c(c2_35_2),.s(s3_36_4),.co(c3_36_4)
);
wire c3_37_1, s3_37_1;
full_adder fa3_37_1 (
.a(s2_37_6),.b(s2_37_5),.c(s2_37_4),.s(s3_37_1),.co(c3_37_1)
);
wire c3_37_2, s3_37_2;
full_adder fa3_37_2 (
.a(s2_37_3),.b(s2_37_2),.c(s2_37_1),.s(s3_37_2),.co(c3_37_2)
);
wire c3_37_3, s3_37_3;
full_adder fa3_37_3 (
.a(c2_36_6),.b(c2_36_5),.c(c2_36_4),.s(s3_37_3),.co(c3_37_3)
);
wire c3_37_4, s3_37_4;
full_adder fa3_37_4 (
.a(c2_36_3),.b(c2_36_2),.c(c2_36_1),.s(s3_37_4),.co(c3_37_4)
);
wire c3_38_1, s3_38_1;
full_adder fa3_38_1 (
.a(s2_38_6),.b(s2_38_5),.c(s2_38_4),.s(s3_38_1),.co(c3_38_1)
);
wire c3_38_2, s3_38_2;
full_adder fa3_38_2 (
.a(s2_38_3),.b(s2_38_2),.c(s2_38_1),.s(s3_38_2),.co(c3_38_2)
);
wire c3_38_3, s3_38_3;
full_adder fa3_38_3 (
.a(c2_37_6),.b(c2_37_5),.c(c2_37_4),.s(s3_38_3),.co(c3_38_3)
);
wire c3_38_4, s3_38_4;
full_adder fa3_38_4 (
.a(c2_37_3),.b(c2_37_2),.c(c2_37_1),.s(s3_38_4),.co(c3_38_4)
);
wire c3_39_1, s3_39_1;
full_adder fa3_39_1 (
.a(c1_38_1),.b(s2_39_5),.c(s2_39_4),.s(s3_39_1),.co(c3_39_1)
);
wire c3_39_2, s3_39_2;
full_adder fa3_39_2 (
.a(s2_39_3),.b(s2_39_2),.c(s2_39_1),.s(s3_39_2),.co(c3_39_2)
);
wire c3_39_3, s3_39_3;
full_adder fa3_39_3 (
.a(c2_38_6),.b(c2_38_5),.c(c2_38_4),.s(s3_39_3),.co(c3_39_3)
);
wire c3_39_4, s3_39_4;
full_adder fa3_39_4 (
.a(c2_38_3),.b(c2_38_2),.c(c2_38_1),.s(s3_39_4),.co(c3_39_4)
);
wire c3_40_1, s3_40_1;
full_adder fa3_40_1 (
.a(c1_39_1),.b(s2_40_5),.c(s2_40_4),.s(s3_40_1),.co(c3_40_1)
);
wire c3_40_2, s3_40_2;
full_adder fa3_40_2 (
.a(s2_40_3),.b(s2_40_2),.c(s2_40_1),.s(s3_40_2),.co(c3_40_2)
);
wire c3_40_3, s3_40_3;
full_adder fa3_40_3 (
.a(c2_39_5),.b(c2_39_4),.c(c2_39_3),.s(s3_40_3),.co(c3_40_3)
);
wire c3_40_4, s3_40_4;
half_adder ha3_40_4 (
.a(c2_39_2),.b(c2_39_1),.p(s3_40_4),.g(c3_40_4)
);
wire c3_41_1, s3_41_1;
full_adder fa3_41_1 (
.a(c1_40_1),.b(s2_41_5),.c(s2_41_4),.s(s3_41_1),.co(c3_41_1)
);
wire c3_41_2, s3_41_2;
full_adder fa3_41_2 (
.a(s2_41_3),.b(s2_41_2),.c(s2_41_1),.s(s3_41_2),.co(c3_41_2)
);
wire c3_41_3, s3_41_3;
full_adder fa3_41_3 (
.a(c2_40_5),.b(c2_40_4),.c(c2_40_3),.s(s3_41_3),.co(c3_41_3)
);
wire c3_41_4, s3_41_4;
half_adder ha3_41_4 (
.a(c2_40_2),.b(c2_40_1),.p(s3_41_4),.g(c3_41_4)
);
wire c3_42_1, s3_42_1;
full_adder fa3_42_1 (
.a(s2_42_5),.b(s2_42_4),.c(s2_42_3),.s(s3_42_1),.co(c3_42_1)
);
wire c3_42_2, s3_42_2;
full_adder fa3_42_2 (
.a(s2_42_2),.b(s2_42_1),.c(c2_41_5),.s(s3_42_2),.co(c3_42_2)
);
wire c3_42_3, s3_42_3;
full_adder fa3_42_3 (
.a(c2_41_4),.b(c2_41_3),.c(c2_41_2),.s(s3_42_3),.co(c3_42_3)
);
wire c3_43_1, s3_43_1;
full_adder fa3_43_1 (
.a(s2_43_5),.b(s2_43_4),.c(s2_43_3),.s(s3_43_1),.co(c3_43_1)
);
wire c3_43_2, s3_43_2;
full_adder fa3_43_2 (
.a(s2_43_2),.b(s2_43_1),.c(c2_42_5),.s(s3_43_2),.co(c3_43_2)
);
wire c3_43_3, s3_43_3;
full_adder fa3_43_3 (
.a(c2_42_4),.b(c2_42_3),.c(c2_42_2),.s(s3_43_3),.co(c3_43_3)
);
wire c3_44_1, s3_44_1;
full_adder fa3_44_1 (
.a(s2_44_5),.b(s2_44_4),.c(s2_44_3),.s(s3_44_1),.co(c3_44_1)
);
wire c3_44_2, s3_44_2;
full_adder fa3_44_2 (
.a(s2_44_2),.b(s2_44_1),.c(c2_43_5),.s(s3_44_2),.co(c3_44_2)
);
wire c3_44_3, s3_44_3;
full_adder fa3_44_3 (
.a(c2_43_4),.b(c2_43_3),.c(c2_43_2),.s(s3_44_3),.co(c3_44_3)
);
wire c3_45_1, s3_45_1;
full_adder fa3_45_1 (
.a(s2_45_4),.b(s2_45_3),.c(s2_45_2),.s(s3_45_1),.co(c3_45_1)
);
wire c3_45_2, s3_45_2;
full_adder fa3_45_2 (
.a(s2_45_1),.b(c2_44_5),.c(c2_44_4),.s(s3_45_2),.co(c3_45_2)
);
wire c3_45_3, s3_45_3;
full_adder fa3_45_3 (
.a(c2_44_3),.b(c2_44_2),.c(c2_44_1),.s(s3_45_3),.co(c3_45_3)
);
wire c3_46_1, s3_46_1;
full_adder fa3_46_1 (
.a(s2_46_4),.b(s2_46_3),.c(s2_46_2),.s(s3_46_1),.co(c3_46_1)
);
wire c3_46_2, s3_46_2;
full_adder fa3_46_2 (
.a(s2_46_1),.b(c2_45_4),.c(c2_45_3),.s(s3_46_2),.co(c3_46_2)
);
wire c3_46_3, s3_46_3;
half_adder ha3_46_3 (
.a(c2_45_2),.b(c2_45_1),.p(s3_46_3),.g(c3_46_3)
);
wire c3_47_1, s3_47_1;
full_adder fa3_47_1 (
.a(s2_47_4),.b(s2_47_3),.c(s2_47_2),.s(s3_47_1),.co(c3_47_1)
);
wire c3_47_2, s3_47_2;
full_adder fa3_47_2 (
.a(s2_47_1),.b(c2_46_4),.c(c2_46_3),.s(s3_47_2),.co(c3_47_2)
);
wire c3_47_3, s3_47_3;
half_adder ha3_47_3 (
.a(c2_46_2),.b(c2_46_1),.p(s3_47_3),.g(c3_47_3)
);
wire c3_48_1, s3_48_1;
full_adder fa3_48_1 (
.a(c1_47_1),.b(s2_48_3),.c(s2_48_2),.s(s3_48_1),.co(c3_48_1)
);
wire c3_48_2, s3_48_2;
full_adder fa3_48_2 (
.a(s2_48_1),.b(c2_47_4),.c(c2_47_3),.s(s3_48_2),.co(c3_48_2)
);
wire c3_48_3, s3_48_3;
half_adder ha3_48_3 (
.a(c2_47_2),.b(c2_47_1),.p(s3_48_3),.g(c3_48_3)
);
wire c3_49_1, s3_49_1;
full_adder fa3_49_1 (
.a(c1_48_1),.b(s2_49_3),.c(s2_49_2),.s(s3_49_1),.co(c3_49_1)
);
wire c3_49_2, s3_49_2;
full_adder fa3_49_2 (
.a(s2_49_1),.b(c2_48_3),.c(c2_48_2),.s(s3_49_2),.co(c3_49_2)
);
wire c3_50_1, s3_50_1;
full_adder fa3_50_1 (
.a(c1_49_1),.b(s2_50_3),.c(s2_50_2),.s(s3_50_1),.co(c3_50_1)
);
wire c3_50_2, s3_50_2;
full_adder fa3_50_2 (
.a(s2_50_1),.b(c2_49_3),.c(c2_49_2),.s(s3_50_2),.co(c3_50_2)
);
wire c3_51_1, s3_51_1;
full_adder fa3_51_1 (
.a(s2_51_3),.b(s2_51_2),.c(s2_51_1),.s(s3_51_1),.co(c3_51_1)
);
wire c3_51_2, s3_51_2;
full_adder fa3_51_2 (
.a(c2_50_3),.b(c2_50_2),.c(c2_50_1),.s(s3_51_2),.co(c3_51_2)
);
wire c3_52_1, s3_52_1;
full_adder fa3_52_1 (
.a(s2_52_3),.b(s2_52_2),.c(s2_52_1),.s(s3_52_1),.co(c3_52_1)
);
wire c3_52_2, s3_52_2;
full_adder fa3_52_2 (
.a(c2_51_3),.b(c2_51_2),.c(c2_51_1),.s(s3_52_2),.co(c3_52_2)
);
wire c3_53_1, s3_53_1;
full_adder fa3_53_1 (
.a(s2_53_3),.b(s2_53_2),.c(s2_53_1),.s(s3_53_1),.co(c3_53_1)
);
wire c3_53_2, s3_53_2;
full_adder fa3_53_2 (
.a(c2_52_3),.b(c2_52_2),.c(c2_52_1),.s(s3_53_2),.co(c3_53_2)
);
wire c3_54_1, s3_54_1;
full_adder fa3_54_1 (
.a(s2_54_2),.b(s2_54_1),.c(c2_53_3),.s(s3_54_1),.co(c3_54_1)
);
wire c3_54_2, s3_54_2;
half_adder ha3_54_2 (
.a(c2_53_2),.b(c2_53_1),.p(s3_54_2),.g(c3_54_2)
);
wire c3_55_1, s3_55_1;
full_adder fa3_55_1 (
.a(s2_55_2),.b(s2_55_1),.c(c2_54_2),.s(s3_55_1),.co(c3_55_1)
);
wire c3_56_1, s3_56_1;
full_adder fa3_56_1 (
.a(s2_56_2),.b(s2_56_1),.c(c2_55_2),.s(s3_56_1),.co(c3_56_1)
);
wire c3_57_1, s3_57_1;
full_adder fa3_57_1 (
.a(c1_56_1),.b(s2_57_1),.c(c2_56_2),.s(s3_57_1),.co(c3_57_1)
);
wire c3_58_1, s3_58_1;
full_adder fa3_58_1 (
.a(c1_57_1),.b(s2_58_1),.c(c2_57_1),.s(s3_58_1),.co(c3_58_1)
);
wire c3_59_1, s3_59_1;
full_adder fa3_59_1 (
.a(c1_58_1),.b(s2_59_1),.c(c2_58_1),.s(s3_59_1),.co(c3_59_1)
);
wire c3_60_1, s3_60_1;
half_adder ha3_60_1 (
.a(s2_60_1),.b(c2_59_1),.p(s3_60_1),.g(c3_60_1)
);
wire c3_61_1, s3_61_1;
half_adder ha3_61_1 (
.a(s2_61_1),.b(c2_60_1),.p(s3_61_1),.g(c3_61_1)
);
wire c3_62_1, s3_62_1;
half_adder ha3_62_1 (
.a(s2_62_1),.b(c2_61_1),.p(s3_62_1),.g(c3_62_1)
);
wire c4_4_1, s4_4_1;
half_adder ha4_4_1 (
.a(s3_4_1),.b(c3_3_1),.p(s4_4_1),.g(c4_4_1)
);
wire c4_5_1, s4_5_1;
half_adder ha4_5_1 (
.a(s3_5_1),.b(c3_4_1),.p(s4_5_1),.g(c4_5_1)
);
wire c4_6_1, s4_6_1;
half_adder ha4_6_1 (
.a(s3_6_1),.b(c3_5_1),.p(s4_6_1),.g(c4_6_1)
);
wire c4_7_1, s4_7_1;
full_adder fa4_7_1 (
.a(c2_6_1),.b(s3_7_1),.c(c3_6_1),.s(s4_7_1),.co(c4_7_1)
);
wire c4_8_1, s4_8_1;
full_adder fa4_8_1 (
.a(c2_7_1),.b(s3_8_1),.c(c3_7_1),.s(s4_8_1),.co(c4_8_1)
);
wire c4_9_1, s4_9_1;
full_adder fa4_9_1 (
.a(s3_9_2),.b(s3_9_1),.c(c3_8_1),.s(s4_9_1),.co(c4_9_1)
);
wire c4_10_1, s4_10_1;
full_adder fa4_10_1 (
.a(s3_10_2),.b(s3_10_1),.c(c3_9_2),.s(s4_10_1),.co(c4_10_1)
);
wire c4_11_1, s4_11_1;
full_adder fa4_11_1 (
.a(s3_11_2),.b(s3_11_1),.c(c3_10_2),.s(s4_11_1),.co(c4_11_1)
);
wire c4_12_1, s4_12_1;
full_adder fa4_12_1 (
.a(s3_12_2),.b(s3_12_1),.c(c3_11_2),.s(s4_12_1),.co(c4_12_1)
);
wire c4_13_1, s4_13_1;
full_adder fa4_13_1 (
.a(s3_13_2),.b(s3_13_1),.c(c3_12_2),.s(s4_13_1),.co(c4_13_1)
);
wire c4_14_1, s4_14_1;
full_adder fa4_14_1 (
.a(c2_13_1),.b(s3_14_2),.c(s3_14_1),.s(s4_14_1),.co(c4_14_1)
);
wire c4_14_2, s4_14_2;
half_adder ha4_14_2 (
.a(c3_13_2),.b(c3_13_1),.p(s4_14_2),.g(c4_14_2)
);
wire c4_15_1, s4_15_1;
full_adder fa4_15_1 (
.a(c2_14_1),.b(s3_15_2),.c(s3_15_1),.s(s4_15_1),.co(c4_15_1)
);
wire c4_15_2, s4_15_2;
half_adder ha4_15_2 (
.a(c3_14_2),.b(c3_14_1),.p(s4_15_2),.g(c4_15_2)
);
wire c4_16_1, s4_16_1;
full_adder fa4_16_1 (
.a(s3_16_3),.b(s3_16_2),.c(s3_16_1),.s(s4_16_1),.co(c4_16_1)
);
wire c4_16_2, s4_16_2;
half_adder ha4_16_2 (
.a(c3_15_2),.b(c3_15_1),.p(s4_16_2),.g(c4_16_2)
);
wire c4_17_1, s4_17_1;
full_adder fa4_17_1 (
.a(s3_17_3),.b(s3_17_2),.c(s3_17_1),.s(s4_17_1),.co(c4_17_1)
);
wire c4_17_2, s4_17_2;
full_adder fa4_17_2 (
.a(c3_16_3),.b(c3_16_2),.c(c3_16_1),.s(s4_17_2),.co(c4_17_2)
);
wire c4_18_1, s4_18_1;
full_adder fa4_18_1 (
.a(s3_18_3),.b(s3_18_2),.c(s3_18_1),.s(s4_18_1),.co(c4_18_1)
);
wire c4_18_2, s4_18_2;
full_adder fa4_18_2 (
.a(c3_17_3),.b(c3_17_2),.c(c3_17_1),.s(s4_18_2),.co(c4_18_2)
);
wire c4_19_1, s4_19_1;
full_adder fa4_19_1 (
.a(s3_19_3),.b(s3_19_2),.c(s3_19_1),.s(s4_19_1),.co(c4_19_1)
);
wire c4_19_2, s4_19_2;
full_adder fa4_19_2 (
.a(c3_18_3),.b(c3_18_2),.c(c3_18_1),.s(s4_19_2),.co(c4_19_2)
);
wire c4_20_1, s4_20_1;
full_adder fa4_20_1 (
.a(s3_20_3),.b(s3_20_2),.c(s3_20_1),.s(s4_20_1),.co(c4_20_1)
);
wire c4_20_2, s4_20_2;
full_adder fa4_20_2 (
.a(c3_19_3),.b(c3_19_2),.c(c3_19_1),.s(s4_20_2),.co(c4_20_2)
);
wire c4_21_1, s4_21_1;
full_adder fa4_21_1 (
.a(c2_20_1),.b(s3_21_3),.c(s3_21_2),.s(s4_21_1),.co(c4_21_1)
);
wire c4_21_2, s4_21_2;
full_adder fa4_21_2 (
.a(s3_21_1),.b(c3_20_3),.c(c3_20_2),.s(s4_21_2),.co(c4_21_2)
);
wire c4_22_1, s4_22_1;
full_adder fa4_22_1 (
.a(c2_21_1),.b(s3_22_3),.c(s3_22_2),.s(s4_22_1),.co(c4_22_1)
);
wire c4_22_2, s4_22_2;
full_adder fa4_22_2 (
.a(s3_22_1),.b(c3_21_3),.c(c3_21_2),.s(s4_22_2),.co(c4_22_2)
);
wire c4_23_1, s4_23_1;
full_adder fa4_23_1 (
.a(s3_23_4),.b(s3_23_3),.c(s3_23_2),.s(s4_23_1),.co(c4_23_1)
);
wire c4_23_2, s4_23_2;
full_adder fa4_23_2 (
.a(s3_23_1),.b(c3_22_3),.c(c3_22_2),.s(s4_23_2),.co(c4_23_2)
);
wire c4_24_1, s4_24_1;
full_adder fa4_24_1 (
.a(s3_24_4),.b(s3_24_3),.c(s3_24_2),.s(s4_24_1),.co(c4_24_1)
);
wire c4_24_2, s4_24_2;
full_adder fa4_24_2 (
.a(s3_24_1),.b(c3_23_4),.c(c3_23_3),.s(s4_24_2),.co(c4_24_2)
);
wire c4_24_3, s4_24_3;
half_adder ha4_24_3 (
.a(c3_23_2),.b(c3_23_1),.p(s4_24_3),.g(c4_24_3)
);
wire c4_25_1, s4_25_1;
full_adder fa4_25_1 (
.a(s3_25_4),.b(s3_25_3),.c(s3_25_2),.s(s4_25_1),.co(c4_25_1)
);
wire c4_25_2, s4_25_2;
full_adder fa4_25_2 (
.a(s3_25_1),.b(c3_24_4),.c(c3_24_3),.s(s4_25_2),.co(c4_25_2)
);
wire c4_25_3, s4_25_3;
half_adder ha4_25_3 (
.a(c3_24_2),.b(c3_24_1),.p(s4_25_3),.g(c4_25_3)
);
wire c4_26_1, s4_26_1;
full_adder fa4_26_1 (
.a(s3_26_4),.b(s3_26_3),.c(s3_26_2),.s(s4_26_1),.co(c4_26_1)
);
wire c4_26_2, s4_26_2;
full_adder fa4_26_2 (
.a(s3_26_1),.b(c3_25_4),.c(c3_25_3),.s(s4_26_2),.co(c4_26_2)
);
wire c4_26_3, s4_26_3;
half_adder ha4_26_3 (
.a(c3_25_2),.b(c3_25_1),.p(s4_26_3),.g(c4_26_3)
);
wire c4_27_1, s4_27_1;
full_adder fa4_27_1 (
.a(c2_26_1),.b(s3_27_4),.c(s3_27_3),.s(s4_27_1),.co(c4_27_1)
);
wire c4_27_2, s4_27_2;
full_adder fa4_27_2 (
.a(s3_27_2),.b(s3_27_1),.c(c3_26_4),.s(s4_27_2),.co(c4_27_2)
);
wire c4_27_3, s4_27_3;
full_adder fa4_27_3 (
.a(c3_26_3),.b(c3_26_2),.c(c3_26_1),.s(s4_27_3),.co(c4_27_3)
);
wire c4_28_1, s4_28_1;
full_adder fa4_28_1 (
.a(c2_27_1),.b(s3_28_4),.c(s3_28_3),.s(s4_28_1),.co(c4_28_1)
);
wire c4_28_2, s4_28_2;
full_adder fa4_28_2 (
.a(s3_28_2),.b(s3_28_1),.c(c3_27_4),.s(s4_28_2),.co(c4_28_2)
);
wire c4_28_3, s4_28_3;
full_adder fa4_28_3 (
.a(c3_27_3),.b(c3_27_2),.c(c3_27_1),.s(s4_28_3),.co(c4_28_3)
);
wire c4_29_1, s4_29_1;
full_adder fa4_29_1 (
.a(c2_28_1),.b(s3_29_4),.c(s3_29_3),.s(s4_29_1),.co(c4_29_1)
);
wire c4_29_2, s4_29_2;
full_adder fa4_29_2 (
.a(s3_29_2),.b(s3_29_1),.c(c3_28_4),.s(s4_29_2),.co(c4_29_2)
);
wire c4_29_3, s4_29_3;
full_adder fa4_29_3 (
.a(c3_28_3),.b(c3_28_2),.c(c3_28_1),.s(s4_29_3),.co(c4_29_3)
);
wire c4_30_1, s4_30_1;
full_adder fa4_30_1 (
.a(s3_30_5),.b(s3_30_4),.c(s3_30_3),.s(s4_30_1),.co(c4_30_1)
);
wire c4_30_2, s4_30_2;
full_adder fa4_30_2 (
.a(s3_30_2),.b(s3_30_1),.c(c3_29_4),.s(s4_30_2),.co(c4_30_2)
);
wire c4_30_3, s4_30_3;
full_adder fa4_30_3 (
.a(c3_29_3),.b(c3_29_2),.c(c3_29_1),.s(s4_30_3),.co(c4_30_3)
);
wire c4_31_1, s4_31_1;
full_adder fa4_31_1 (
.a(s3_31_5),.b(s3_31_4),.c(s3_31_3),.s(s4_31_1),.co(c4_31_1)
);
wire c4_31_2, s4_31_2;
full_adder fa4_31_2 (
.a(s3_31_2),.b(s3_31_1),.c(c3_30_5),.s(s4_31_2),.co(c4_31_2)
);
wire c4_31_3, s4_31_3;
full_adder fa4_31_3 (
.a(c3_30_4),.b(c3_30_3),.c(c3_30_2),.s(s4_31_3),.co(c4_31_3)
);
wire c4_32_1, s4_32_1;
full_adder fa4_32_1 (
.a(s3_32_5),.b(s3_32_4),.c(s3_32_3),.s(s4_32_1),.co(c4_32_1)
);
wire c4_32_2, s4_32_2;
full_adder fa4_32_2 (
.a(s3_32_2),.b(s3_32_1),.c(c3_31_5),.s(s4_32_2),.co(c4_32_2)
);
wire c4_32_3, s4_32_3;
full_adder fa4_32_3 (
.a(c3_31_4),.b(c3_31_3),.c(c3_31_2),.s(s4_32_3),.co(c4_32_3)
);
wire c4_33_1, s4_33_1;
full_adder fa4_33_1 (
.a(s3_33_5),.b(s3_33_4),.c(s3_33_3),.s(s4_33_1),.co(c4_33_1)
);
wire c4_33_2, s4_33_2;
full_adder fa4_33_2 (
.a(s3_33_2),.b(s3_33_1),.c(c3_32_5),.s(s4_33_2),.co(c4_33_2)
);
wire c4_33_3, s4_33_3;
full_adder fa4_33_3 (
.a(c3_32_4),.b(c3_32_3),.c(c3_32_2),.s(s4_33_3),.co(c4_33_3)
);
wire c4_34_1, s4_34_1;
full_adder fa4_34_1 (
.a(s3_34_5),.b(s3_34_4),.c(s3_34_3),.s(s4_34_1),.co(c4_34_1)
);
wire c4_34_2, s4_34_2;
full_adder fa4_34_2 (
.a(s3_34_2),.b(s3_34_1),.c(c3_33_5),.s(s4_34_2),.co(c4_34_2)
);
wire c4_34_3, s4_34_3;
full_adder fa4_34_3 (
.a(c3_33_4),.b(c3_33_3),.c(c3_33_2),.s(s4_34_3),.co(c4_34_3)
);
wire c4_35_1, s4_35_1;
full_adder fa4_35_1 (
.a(s3_35_5),.b(s3_35_4),.c(s3_35_3),.s(s4_35_1),.co(c4_35_1)
);
wire c4_35_2, s4_35_2;
full_adder fa4_35_2 (
.a(s3_35_2),.b(s3_35_1),.c(c3_34_5),.s(s4_35_2),.co(c4_35_2)
);
wire c4_35_3, s4_35_3;
full_adder fa4_35_3 (
.a(c3_34_4),.b(c3_34_3),.c(c3_34_2),.s(s4_35_3),.co(c4_35_3)
);
wire c4_36_1, s4_36_1;
full_adder fa4_36_1 (
.a(c2_35_1),.b(s3_36_4),.c(s3_36_3),.s(s4_36_1),.co(c4_36_1)
);
wire c4_36_2, s4_36_2;
full_adder fa4_36_2 (
.a(s3_36_2),.b(s3_36_1),.c(c3_35_5),.s(s4_36_2),.co(c4_36_2)
);
wire c4_36_3, s4_36_3;
full_adder fa4_36_3 (
.a(c3_35_4),.b(c3_35_3),.c(c3_35_2),.s(s4_36_3),.co(c4_36_3)
);
wire c4_37_1, s4_37_1;
full_adder fa4_37_1 (
.a(s3_37_4),.b(s3_37_3),.c(s3_37_2),.s(s4_37_1),.co(c4_37_1)
);
wire c4_37_2, s4_37_2;
full_adder fa4_37_2 (
.a(s3_37_1),.b(c3_36_4),.c(c3_36_3),.s(s4_37_2),.co(c4_37_2)
);
wire c4_37_3, s4_37_3;
half_adder ha4_37_3 (
.a(c3_36_2),.b(c3_36_1),.p(s4_37_3),.g(c4_37_3)
);
wire c4_38_1, s4_38_1;
full_adder fa4_38_1 (
.a(s3_38_4),.b(s3_38_3),.c(s3_38_2),.s(s4_38_1),.co(c4_38_1)
);
wire c4_38_2, s4_38_2;
full_adder fa4_38_2 (
.a(s3_38_1),.b(c3_37_4),.c(c3_37_3),.s(s4_38_2),.co(c4_38_2)
);
wire c4_38_3, s4_38_3;
half_adder ha4_38_3 (
.a(c3_37_2),.b(c3_37_1),.p(s4_38_3),.g(c4_38_3)
);
wire c4_39_1, s4_39_1;
full_adder fa4_39_1 (
.a(s3_39_4),.b(s3_39_3),.c(s3_39_2),.s(s4_39_1),.co(c4_39_1)
);
wire c4_39_2, s4_39_2;
full_adder fa4_39_2 (
.a(s3_39_1),.b(c3_38_4),.c(c3_38_3),.s(s4_39_2),.co(c4_39_2)
);
wire c4_39_3, s4_39_3;
half_adder ha4_39_3 (
.a(c3_38_2),.b(c3_38_1),.p(s4_39_3),.g(c4_39_3)
);
wire c4_40_1, s4_40_1;
full_adder fa4_40_1 (
.a(s3_40_4),.b(s3_40_3),.c(s3_40_2),.s(s4_40_1),.co(c4_40_1)
);
wire c4_40_2, s4_40_2;
full_adder fa4_40_2 (
.a(s3_40_1),.b(c3_39_4),.c(c3_39_3),.s(s4_40_2),.co(c4_40_2)
);
wire c4_40_3, s4_40_3;
half_adder ha4_40_3 (
.a(c3_39_2),.b(c3_39_1),.p(s4_40_3),.g(c4_40_3)
);
wire c4_41_1, s4_41_1;
full_adder fa4_41_1 (
.a(s3_41_4),.b(s3_41_3),.c(s3_41_2),.s(s4_41_1),.co(c4_41_1)
);
wire c4_41_2, s4_41_2;
full_adder fa4_41_2 (
.a(s3_41_1),.b(c3_40_4),.c(c3_40_3),.s(s4_41_2),.co(c4_41_2)
);
wire c4_41_3, s4_41_3;
half_adder ha4_41_3 (
.a(c3_40_2),.b(c3_40_1),.p(s4_41_3),.g(c4_41_3)
);
wire c4_42_1, s4_42_1;
full_adder fa4_42_1 (
.a(c2_41_1),.b(s3_42_3),.c(s3_42_2),.s(s4_42_1),.co(c4_42_1)
);
wire c4_42_2, s4_42_2;
full_adder fa4_42_2 (
.a(s3_42_1),.b(c3_41_4),.c(c3_41_3),.s(s4_42_2),.co(c4_42_2)
);
wire c4_42_3, s4_42_3;
half_adder ha4_42_3 (
.a(c3_41_2),.b(c3_41_1),.p(s4_42_3),.g(c4_42_3)
);
wire c4_43_1, s4_43_1;
full_adder fa4_43_1 (
.a(c2_42_1),.b(s3_43_3),.c(s3_43_2),.s(s4_43_1),.co(c4_43_1)
);
wire c4_43_2, s4_43_2;
full_adder fa4_43_2 (
.a(s3_43_1),.b(c3_42_3),.c(c3_42_2),.s(s4_43_2),.co(c4_43_2)
);
wire c4_44_1, s4_44_1;
full_adder fa4_44_1 (
.a(c2_43_1),.b(s3_44_3),.c(s3_44_2),.s(s4_44_1),.co(c4_44_1)
);
wire c4_44_2, s4_44_2;
full_adder fa4_44_2 (
.a(s3_44_1),.b(c3_43_3),.c(c3_43_2),.s(s4_44_2),.co(c4_44_2)
);
wire c4_45_1, s4_45_1;
full_adder fa4_45_1 (
.a(s3_45_3),.b(s3_45_2),.c(s3_45_1),.s(s4_45_1),.co(c4_45_1)
);
wire c4_45_2, s4_45_2;
full_adder fa4_45_2 (
.a(c3_44_3),.b(c3_44_2),.c(c3_44_1),.s(s4_45_2),.co(c4_45_2)
);
wire c4_46_1, s4_46_1;
full_adder fa4_46_1 (
.a(s3_46_3),.b(s3_46_2),.c(s3_46_1),.s(s4_46_1),.co(c4_46_1)
);
wire c4_46_2, s4_46_2;
full_adder fa4_46_2 (
.a(c3_45_3),.b(c3_45_2),.c(c3_45_1),.s(s4_46_2),.co(c4_46_2)
);
wire c4_47_1, s4_47_1;
full_adder fa4_47_1 (
.a(s3_47_3),.b(s3_47_2),.c(s3_47_1),.s(s4_47_1),.co(c4_47_1)
);
wire c4_47_2, s4_47_2;
full_adder fa4_47_2 (
.a(c3_46_3),.b(c3_46_2),.c(c3_46_1),.s(s4_47_2),.co(c4_47_2)
);
wire c4_48_1, s4_48_1;
full_adder fa4_48_1 (
.a(s3_48_3),.b(s3_48_2),.c(s3_48_1),.s(s4_48_1),.co(c4_48_1)
);
wire c4_48_2, s4_48_2;
full_adder fa4_48_2 (
.a(c3_47_3),.b(c3_47_2),.c(c3_47_1),.s(s4_48_2),.co(c4_48_2)
);
wire c4_49_1, s4_49_1;
full_adder fa4_49_1 (
.a(c2_48_1),.b(s3_49_2),.c(s3_49_1),.s(s4_49_1),.co(c4_49_1)
);
wire c4_49_2, s4_49_2;
full_adder fa4_49_2 (
.a(c3_48_3),.b(c3_48_2),.c(c3_48_1),.s(s4_49_2),.co(c4_49_2)
);
wire c4_50_1, s4_50_1;
full_adder fa4_50_1 (
.a(c2_49_1),.b(s3_50_2),.c(s3_50_1),.s(s4_50_1),.co(c4_50_1)
);
wire c4_50_2, s4_50_2;
half_adder ha4_50_2 (
.a(c3_49_2),.b(c3_49_1),.p(s4_50_2),.g(c4_50_2)
);
wire c4_51_1, s4_51_1;
full_adder fa4_51_1 (
.a(s3_51_2),.b(s3_51_1),.c(c3_50_2),.s(s4_51_1),.co(c4_51_1)
);
wire c4_52_1, s4_52_1;
full_adder fa4_52_1 (
.a(s3_52_2),.b(s3_52_1),.c(c3_51_2),.s(s4_52_1),.co(c4_52_1)
);
wire c4_53_1, s4_53_1;
full_adder fa4_53_1 (
.a(s3_53_2),.b(s3_53_1),.c(c3_52_2),.s(s4_53_1),.co(c4_53_1)
);
wire c4_54_1, s4_54_1;
full_adder fa4_54_1 (
.a(s3_54_2),.b(s3_54_1),.c(c3_53_2),.s(s4_54_1),.co(c4_54_1)
);
wire c4_55_1, s4_55_1;
full_adder fa4_55_1 (
.a(c2_54_1),.b(s3_55_1),.c(c3_54_2),.s(s4_55_1),.co(c4_55_1)
);
wire c4_56_1, s4_56_1;
full_adder fa4_56_1 (
.a(c2_55_1),.b(s3_56_1),.c(c3_55_1),.s(s4_56_1),.co(c4_56_1)
);
wire c4_57_1, s4_57_1;
full_adder fa4_57_1 (
.a(c2_56_1),.b(s3_57_1),.c(c3_56_1),.s(s4_57_1),.co(c4_57_1)
);
wire c4_58_1, s4_58_1;
half_adder ha4_58_1 (
.a(s3_58_1),.b(c3_57_1),.p(s4_58_1),.g(c4_58_1)
);
wire c4_59_1, s4_59_1;
half_adder ha4_59_1 (
.a(s3_59_1),.b(c3_58_1),.p(s4_59_1),.g(c4_59_1)
);
wire c4_60_1, s4_60_1;
half_adder ha4_60_1 (
.a(s3_60_1),.b(c3_59_1),.p(s4_60_1),.g(c4_60_1)
);
wire c4_61_1, s4_61_1;
half_adder ha4_61_1 (
.a(s3_61_1),.b(c3_60_1),.p(s4_61_1),.g(c4_61_1)
);
wire c4_62_1, s4_62_1;
half_adder ha4_62_1 (
.a(s3_62_1),.b(c3_61_1),.p(s4_62_1),.g(c4_62_1)
);
wire c4_63_1, s4_63_1;
half_adder ha4_63_1 (
.a(c2_62_1),.b(c3_62_1),.p(s4_63_1),.g(c4_63_1)
);
wire c5_5_1, s5_5_1;
half_adder ha5_5_1 (
.a(s4_5_1),.b(c4_4_1),.p(s5_5_1),.g(c5_5_1)
);
wire c5_6_1, s5_6_1;
half_adder ha5_6_1 (
.a(s4_6_1),.b(c4_5_1),.p(s5_6_1),.g(c5_6_1)
);
wire c5_7_1, s5_7_1;
half_adder ha5_7_1 (
.a(s4_7_1),.b(c4_6_1),.p(s5_7_1),.g(c5_7_1)
);
wire c5_8_1, s5_8_1;
half_adder ha5_8_1 (
.a(s4_8_1),.b(c4_7_1),.p(s5_8_1),.g(c5_8_1)
);
wire c5_9_1, s5_9_1;
half_adder ha5_9_1 (
.a(s4_9_1),.b(c4_8_1),.p(s5_9_1),.g(c5_9_1)
);
wire c5_10_1, s5_10_1;
full_adder fa5_10_1 (
.a(c3_9_1),.b(s4_10_1),.c(c4_9_1),.s(s5_10_1),.co(c5_10_1)
);
wire c5_11_1, s5_11_1;
full_adder fa5_11_1 (
.a(c3_10_1),.b(s4_11_1),.c(c4_10_1),.s(s5_11_1),.co(c5_11_1)
);
wire c5_12_1, s5_12_1;
full_adder fa5_12_1 (
.a(c3_11_1),.b(s4_12_1),.c(c4_11_1),.s(s5_12_1),.co(c5_12_1)
);
wire c5_13_1, s5_13_1;
full_adder fa5_13_1 (
.a(c3_12_1),.b(s4_13_1),.c(c4_12_1),.s(s5_13_1),.co(c5_13_1)
);
wire c5_14_1, s5_14_1;
full_adder fa5_14_1 (
.a(s4_14_2),.b(s4_14_1),.c(c4_13_1),.s(s5_14_1),.co(c5_14_1)
);
wire c5_15_1, s5_15_1;
full_adder fa5_15_1 (
.a(s4_15_2),.b(s4_15_1),.c(c4_14_2),.s(s5_15_1),.co(c5_15_1)
);
wire c5_16_1, s5_16_1;
full_adder fa5_16_1 (
.a(s4_16_2),.b(s4_16_1),.c(c4_15_2),.s(s5_16_1),.co(c5_16_1)
);
wire c5_17_1, s5_17_1;
full_adder fa5_17_1 (
.a(s4_17_2),.b(s4_17_1),.c(c4_16_2),.s(s5_17_1),.co(c5_17_1)
);
wire c5_18_1, s5_18_1;
full_adder fa5_18_1 (
.a(s4_18_2),.b(s4_18_1),.c(c4_17_2),.s(s5_18_1),.co(c5_18_1)
);
wire c5_19_1, s5_19_1;
full_adder fa5_19_1 (
.a(s4_19_2),.b(s4_19_1),.c(c4_18_2),.s(s5_19_1),.co(c5_19_1)
);
wire c5_20_1, s5_20_1;
full_adder fa5_20_1 (
.a(s4_20_2),.b(s4_20_1),.c(c4_19_2),.s(s5_20_1),.co(c5_20_1)
);
wire c5_21_1, s5_21_1;
full_adder fa5_21_1 (
.a(c3_20_1),.b(s4_21_2),.c(s4_21_1),.s(s5_21_1),.co(c5_21_1)
);
wire c5_21_2, s5_21_2;
half_adder ha5_21_2 (
.a(c4_20_2),.b(c4_20_1),.p(s5_21_2),.g(c5_21_2)
);
wire c5_22_1, s5_22_1;
full_adder fa5_22_1 (
.a(c3_21_1),.b(s4_22_2),.c(s4_22_1),.s(s5_22_1),.co(c5_22_1)
);
wire c5_22_2, s5_22_2;
half_adder ha5_22_2 (
.a(c4_21_2),.b(c4_21_1),.p(s5_22_2),.g(c5_22_2)
);
wire c5_23_1, s5_23_1;
full_adder fa5_23_1 (
.a(c3_22_1),.b(s4_23_2),.c(s4_23_1),.s(s5_23_1),.co(c5_23_1)
);
wire c5_23_2, s5_23_2;
half_adder ha5_23_2 (
.a(c4_22_2),.b(c4_22_1),.p(s5_23_2),.g(c5_23_2)
);
wire c5_24_1, s5_24_1;
full_adder fa5_24_1 (
.a(s4_24_3),.b(s4_24_2),.c(s4_24_1),.s(s5_24_1),.co(c5_24_1)
);
wire c5_24_2, s5_24_2;
half_adder ha5_24_2 (
.a(c4_23_2),.b(c4_23_1),.p(s5_24_2),.g(c5_24_2)
);
wire c5_25_1, s5_25_1;
full_adder fa5_25_1 (
.a(s4_25_3),.b(s4_25_2),.c(s4_25_1),.s(s5_25_1),.co(c5_25_1)
);
wire c5_25_2, s5_25_2;
full_adder fa5_25_2 (
.a(c4_24_3),.b(c4_24_2),.c(c4_24_1),.s(s5_25_2),.co(c5_25_2)
);
wire c5_26_1, s5_26_1;
full_adder fa5_26_1 (
.a(s4_26_3),.b(s4_26_2),.c(s4_26_1),.s(s5_26_1),.co(c5_26_1)
);
wire c5_26_2, s5_26_2;
full_adder fa5_26_2 (
.a(c4_25_3),.b(c4_25_2),.c(c4_25_1),.s(s5_26_2),.co(c5_26_2)
);
wire c5_27_1, s5_27_1;
full_adder fa5_27_1 (
.a(s4_27_3),.b(s4_27_2),.c(s4_27_1),.s(s5_27_1),.co(c5_27_1)
);
wire c5_27_2, s5_27_2;
full_adder fa5_27_2 (
.a(c4_26_3),.b(c4_26_2),.c(c4_26_1),.s(s5_27_2),.co(c5_27_2)
);
wire c5_28_1, s5_28_1;
full_adder fa5_28_1 (
.a(s4_28_3),.b(s4_28_2),.c(s4_28_1),.s(s5_28_1),.co(c5_28_1)
);
wire c5_28_2, s5_28_2;
full_adder fa5_28_2 (
.a(c4_27_3),.b(c4_27_2),.c(c4_27_1),.s(s5_28_2),.co(c5_28_2)
);
wire c5_29_1, s5_29_1;
full_adder fa5_29_1 (
.a(s4_29_3),.b(s4_29_2),.c(s4_29_1),.s(s5_29_1),.co(c5_29_1)
);
wire c5_29_2, s5_29_2;
full_adder fa5_29_2 (
.a(c4_28_3),.b(c4_28_2),.c(c4_28_1),.s(s5_29_2),.co(c5_29_2)
);
wire c5_30_1, s5_30_1;
full_adder fa5_30_1 (
.a(s4_30_3),.b(s4_30_2),.c(s4_30_1),.s(s5_30_1),.co(c5_30_1)
);
wire c5_30_2, s5_30_2;
full_adder fa5_30_2 (
.a(c4_29_3),.b(c4_29_2),.c(c4_29_1),.s(s5_30_2),.co(c5_30_2)
);
wire c5_31_1, s5_31_1;
full_adder fa5_31_1 (
.a(c3_30_1),.b(s4_31_3),.c(s4_31_2),.s(s5_31_1),.co(c5_31_1)
);
wire c5_31_2, s5_31_2;
full_adder fa5_31_2 (
.a(s4_31_1),.b(c4_30_3),.c(c4_30_2),.s(s5_31_2),.co(c5_31_2)
);
wire c5_32_1, s5_32_1;
full_adder fa5_32_1 (
.a(c3_31_1),.b(s4_32_3),.c(s4_32_2),.s(s5_32_1),.co(c5_32_1)
);
wire c5_32_2, s5_32_2;
full_adder fa5_32_2 (
.a(s4_32_1),.b(c4_31_3),.c(c4_31_2),.s(s5_32_2),.co(c5_32_2)
);
wire c5_33_1, s5_33_1;
full_adder fa5_33_1 (
.a(c3_32_1),.b(s4_33_3),.c(s4_33_2),.s(s5_33_1),.co(c5_33_1)
);
wire c5_33_2, s5_33_2;
full_adder fa5_33_2 (
.a(s4_33_1),.b(c4_32_3),.c(c4_32_2),.s(s5_33_2),.co(c5_33_2)
);
wire c5_34_1, s5_34_1;
full_adder fa5_34_1 (
.a(c3_33_1),.b(s4_34_3),.c(s4_34_2),.s(s5_34_1),.co(c5_34_1)
);
wire c5_34_2, s5_34_2;
full_adder fa5_34_2 (
.a(s4_34_1),.b(c4_33_3),.c(c4_33_2),.s(s5_34_2),.co(c5_34_2)
);
wire c5_35_1, s5_35_1;
full_adder fa5_35_1 (
.a(c3_34_1),.b(s4_35_3),.c(s4_35_2),.s(s5_35_1),.co(c5_35_1)
);
wire c5_35_2, s5_35_2;
full_adder fa5_35_2 (
.a(s4_35_1),.b(c4_34_3),.c(c4_34_2),.s(s5_35_2),.co(c5_35_2)
);
wire c5_36_1, s5_36_1;
full_adder fa5_36_1 (
.a(c3_35_1),.b(s4_36_3),.c(s4_36_2),.s(s5_36_1),.co(c5_36_1)
);
wire c5_36_2, s5_36_2;
full_adder fa5_36_2 (
.a(s4_36_1),.b(c4_35_3),.c(c4_35_2),.s(s5_36_2),.co(c5_36_2)
);
wire c5_37_1, s5_37_1;
full_adder fa5_37_1 (
.a(s4_37_3),.b(s4_37_2),.c(s4_37_1),.s(s5_37_1),.co(c5_37_1)
);
wire c5_37_2, s5_37_2;
full_adder fa5_37_2 (
.a(c4_36_3),.b(c4_36_2),.c(c4_36_1),.s(s5_37_2),.co(c5_37_2)
);
wire c5_38_1, s5_38_1;
full_adder fa5_38_1 (
.a(s4_38_3),.b(s4_38_2),.c(s4_38_1),.s(s5_38_1),.co(c5_38_1)
);
wire c5_38_2, s5_38_2;
full_adder fa5_38_2 (
.a(c4_37_3),.b(c4_37_2),.c(c4_37_1),.s(s5_38_2),.co(c5_38_2)
);
wire c5_39_1, s5_39_1;
full_adder fa5_39_1 (
.a(s4_39_3),.b(s4_39_2),.c(s4_39_1),.s(s5_39_1),.co(c5_39_1)
);
wire c5_39_2, s5_39_2;
full_adder fa5_39_2 (
.a(c4_38_3),.b(c4_38_2),.c(c4_38_1),.s(s5_39_2),.co(c5_39_2)
);
wire c5_40_1, s5_40_1;
full_adder fa5_40_1 (
.a(s4_40_3),.b(s4_40_2),.c(s4_40_1),.s(s5_40_1),.co(c5_40_1)
);
wire c5_40_2, s5_40_2;
full_adder fa5_40_2 (
.a(c4_39_3),.b(c4_39_2),.c(c4_39_1),.s(s5_40_2),.co(c5_40_2)
);
wire c5_41_1, s5_41_1;
full_adder fa5_41_1 (
.a(s4_41_3),.b(s4_41_2),.c(s4_41_1),.s(s5_41_1),.co(c5_41_1)
);
wire c5_41_2, s5_41_2;
full_adder fa5_41_2 (
.a(c4_40_3),.b(c4_40_2),.c(c4_40_1),.s(s5_41_2),.co(c5_41_2)
);
wire c5_42_1, s5_42_1;
full_adder fa5_42_1 (
.a(s4_42_3),.b(s4_42_2),.c(s4_42_1),.s(s5_42_1),.co(c5_42_1)
);
wire c5_42_2, s5_42_2;
full_adder fa5_42_2 (
.a(c4_41_3),.b(c4_41_2),.c(c4_41_1),.s(s5_42_2),.co(c5_42_2)
);
wire c5_43_1, s5_43_1;
full_adder fa5_43_1 (
.a(c3_42_1),.b(s4_43_2),.c(s4_43_1),.s(s5_43_1),.co(c5_43_1)
);
wire c5_43_2, s5_43_2;
full_adder fa5_43_2 (
.a(c4_42_3),.b(c4_42_2),.c(c4_42_1),.s(s5_43_2),.co(c5_43_2)
);
wire c5_44_1, s5_44_1;
full_adder fa5_44_1 (
.a(c3_43_1),.b(s4_44_2),.c(s4_44_1),.s(s5_44_1),.co(c5_44_1)
);
wire c5_44_2, s5_44_2;
half_adder ha5_44_2 (
.a(c4_43_2),.b(c4_43_1),.p(s5_44_2),.g(c5_44_2)
);
wire c5_45_1, s5_45_1;
full_adder fa5_45_1 (
.a(s4_45_2),.b(s4_45_1),.c(c4_44_2),.s(s5_45_1),.co(c5_45_1)
);
wire c5_46_1, s5_46_1;
full_adder fa5_46_1 (
.a(s4_46_2),.b(s4_46_1),.c(c4_45_2),.s(s5_46_1),.co(c5_46_1)
);
wire c5_47_1, s5_47_1;
full_adder fa5_47_1 (
.a(s4_47_2),.b(s4_47_1),.c(c4_46_2),.s(s5_47_1),.co(c5_47_1)
);
wire c5_48_1, s5_48_1;
full_adder fa5_48_1 (
.a(s4_48_2),.b(s4_48_1),.c(c4_47_2),.s(s5_48_1),.co(c5_48_1)
);
wire c5_49_1, s5_49_1;
full_adder fa5_49_1 (
.a(s4_49_2),.b(s4_49_1),.c(c4_48_2),.s(s5_49_1),.co(c5_49_1)
);
wire c5_50_1, s5_50_1;
full_adder fa5_50_1 (
.a(s4_50_2),.b(s4_50_1),.c(c4_49_2),.s(s5_50_1),.co(c5_50_1)
);
wire c5_51_1, s5_51_1;
full_adder fa5_51_1 (
.a(c3_50_1),.b(s4_51_1),.c(c4_50_2),.s(s5_51_1),.co(c5_51_1)
);
wire c5_52_1, s5_52_1;
full_adder fa5_52_1 (
.a(c3_51_1),.b(s4_52_1),.c(c4_51_1),.s(s5_52_1),.co(c5_52_1)
);
wire c5_53_1, s5_53_1;
full_adder fa5_53_1 (
.a(c3_52_1),.b(s4_53_1),.c(c4_52_1),.s(s5_53_1),.co(c5_53_1)
);
wire c5_54_1, s5_54_1;
full_adder fa5_54_1 (
.a(c3_53_1),.b(s4_54_1),.c(c4_53_1),.s(s5_54_1),.co(c5_54_1)
);
wire c5_55_1, s5_55_1;
full_adder fa5_55_1 (
.a(c3_54_1),.b(s4_55_1),.c(c4_54_1),.s(s5_55_1),.co(c5_55_1)
);
wire c5_56_1, s5_56_1;
half_adder ha5_56_1 (
.a(s4_56_1),.b(c4_55_1),.p(s5_56_1),.g(c5_56_1)
);
wire c5_57_1, s5_57_1;
half_adder ha5_57_1 (
.a(s4_57_1),.b(c4_56_1),.p(s5_57_1),.g(c5_57_1)
);
wire c5_58_1, s5_58_1;
half_adder ha5_58_1 (
.a(s4_58_1),.b(c4_57_1),.p(s5_58_1),.g(c5_58_1)
);
wire c5_59_1, s5_59_1;
half_adder ha5_59_1 (
.a(s4_59_1),.b(c4_58_1),.p(s5_59_1),.g(c5_59_1)
);
wire c5_60_1, s5_60_1;
half_adder ha5_60_1 (
.a(s4_60_1),.b(c4_59_1),.p(s5_60_1),.g(c5_60_1)
);
wire c5_61_1, s5_61_1;
half_adder ha5_61_1 (
.a(s4_61_1),.b(c4_60_1),.p(s5_61_1),.g(c5_61_1)
);
wire c5_62_1, s5_62_1;
half_adder ha5_62_1 (
.a(s4_62_1),.b(c4_61_1),.p(s5_62_1),.g(c5_62_1)
);
wire c5_63_1, s5_63_1;
half_adder ha5_63_1 (
.a(s4_63_1),.b(c4_62_1),.p(s5_63_1),.g(c5_63_1)
);
wire c6_6_1, s6_6_1;
half_adder ha6_6_1 (
.a(s5_6_1),.b(c5_5_1),.p(s6_6_1),.g(c6_6_1)
);
wire c6_7_1, s6_7_1;
half_adder ha6_7_1 (
.a(s5_7_1),.b(c5_6_1),.p(s6_7_1),.g(c6_7_1)
);
wire c6_8_1, s6_8_1;
half_adder ha6_8_1 (
.a(s5_8_1),.b(c5_7_1),.p(s6_8_1),.g(c6_8_1)
);
wire c6_9_1, s6_9_1;
half_adder ha6_9_1 (
.a(s5_9_1),.b(c5_8_1),.p(s6_9_1),.g(c6_9_1)
);
wire c6_10_1, s6_10_1;
half_adder ha6_10_1 (
.a(s5_10_1),.b(c5_9_1),.p(s6_10_1),.g(c6_10_1)
);
wire c6_11_1, s6_11_1;
half_adder ha6_11_1 (
.a(s5_11_1),.b(c5_10_1),.p(s6_11_1),.g(c6_11_1)
);
wire c6_12_1, s6_12_1;
half_adder ha6_12_1 (
.a(s5_12_1),.b(c5_11_1),.p(s6_12_1),.g(c6_12_1)
);
wire c6_13_1, s6_13_1;
half_adder ha6_13_1 (
.a(s5_13_1),.b(c5_12_1),.p(s6_13_1),.g(c6_13_1)
);
wire c6_14_1, s6_14_1;
half_adder ha6_14_1 (
.a(s5_14_1),.b(c5_13_1),.p(s6_14_1),.g(c6_14_1)
);
wire c6_15_1, s6_15_1;
full_adder fa6_15_1 (
.a(c4_14_1),.b(s5_15_1),.c(c5_14_1),.s(s6_15_1),.co(c6_15_1)
);
wire c6_16_1, s6_16_1;
full_adder fa6_16_1 (
.a(c4_15_1),.b(s5_16_1),.c(c5_15_1),.s(s6_16_1),.co(c6_16_1)
);
wire c6_17_1, s6_17_1;
full_adder fa6_17_1 (
.a(c4_16_1),.b(s5_17_1),.c(c5_16_1),.s(s6_17_1),.co(c6_17_1)
);
wire c6_18_1, s6_18_1;
full_adder fa6_18_1 (
.a(c4_17_1),.b(s5_18_1),.c(c5_17_1),.s(s6_18_1),.co(c6_18_1)
);
wire c6_19_1, s6_19_1;
full_adder fa6_19_1 (
.a(c4_18_1),.b(s5_19_1),.c(c5_18_1),.s(s6_19_1),.co(c6_19_1)
);
wire c6_20_1, s6_20_1;
full_adder fa6_20_1 (
.a(c4_19_1),.b(s5_20_1),.c(c5_19_1),.s(s6_20_1),.co(c6_20_1)
);
wire c6_21_1, s6_21_1;
full_adder fa6_21_1 (
.a(s5_21_2),.b(s5_21_1),.c(c5_20_1),.s(s6_21_1),.co(c6_21_1)
);
wire c6_22_1, s6_22_1;
full_adder fa6_22_1 (
.a(s5_22_2),.b(s5_22_1),.c(c5_21_2),.s(s6_22_1),.co(c6_22_1)
);
wire c6_23_1, s6_23_1;
full_adder fa6_23_1 (
.a(s5_23_2),.b(s5_23_1),.c(c5_22_2),.s(s6_23_1),.co(c6_23_1)
);
wire c6_24_1, s6_24_1;
full_adder fa6_24_1 (
.a(s5_24_2),.b(s5_24_1),.c(c5_23_2),.s(s6_24_1),.co(c6_24_1)
);
wire c6_25_1, s6_25_1;
full_adder fa6_25_1 (
.a(s5_25_2),.b(s5_25_1),.c(c5_24_2),.s(s6_25_1),.co(c6_25_1)
);
wire c6_26_1, s6_26_1;
full_adder fa6_26_1 (
.a(s5_26_2),.b(s5_26_1),.c(c5_25_2),.s(s6_26_1),.co(c6_26_1)
);
wire c6_27_1, s6_27_1;
full_adder fa6_27_1 (
.a(s5_27_2),.b(s5_27_1),.c(c5_26_2),.s(s6_27_1),.co(c6_27_1)
);
wire c6_28_1, s6_28_1;
full_adder fa6_28_1 (
.a(s5_28_2),.b(s5_28_1),.c(c5_27_2),.s(s6_28_1),.co(c6_28_1)
);
wire c6_29_1, s6_29_1;
full_adder fa6_29_1 (
.a(s5_29_2),.b(s5_29_1),.c(c5_28_2),.s(s6_29_1),.co(c6_29_1)
);
wire c6_30_1, s6_30_1;
full_adder fa6_30_1 (
.a(s5_30_2),.b(s5_30_1),.c(c5_29_2),.s(s6_30_1),.co(c6_30_1)
);
wire c6_31_1, s6_31_1;
full_adder fa6_31_1 (
.a(c4_30_1),.b(s5_31_2),.c(s5_31_1),.s(s6_31_1),.co(c6_31_1)
);
wire c6_31_2, s6_31_2;
half_adder ha6_31_2 (
.a(c5_30_2),.b(c5_30_1),.p(s6_31_2),.g(c6_31_2)
);
wire c6_32_1, s6_32_1;
full_adder fa6_32_1 (
.a(c4_31_1),.b(s5_32_2),.c(s5_32_1),.s(s6_32_1),.co(c6_32_1)
);
wire c6_32_2, s6_32_2;
half_adder ha6_32_2 (
.a(c5_31_2),.b(c5_31_1),.p(s6_32_2),.g(c6_32_2)
);
wire c6_33_1, s6_33_1;
full_adder fa6_33_1 (
.a(c4_32_1),.b(s5_33_2),.c(s5_33_1),.s(s6_33_1),.co(c6_33_1)
);
wire c6_33_2, s6_33_2;
half_adder ha6_33_2 (
.a(c5_32_2),.b(c5_32_1),.p(s6_33_2),.g(c6_33_2)
);
wire c6_34_1, s6_34_1;
full_adder fa6_34_1 (
.a(c4_33_1),.b(s5_34_2),.c(s5_34_1),.s(s6_34_1),.co(c6_34_1)
);
wire c6_34_2, s6_34_2;
half_adder ha6_34_2 (
.a(c5_33_2),.b(c5_33_1),.p(s6_34_2),.g(c6_34_2)
);
wire c6_35_1, s6_35_1;
full_adder fa6_35_1 (
.a(c4_34_1),.b(s5_35_2),.c(s5_35_1),.s(s6_35_1),.co(c6_35_1)
);
wire c6_35_2, s6_35_2;
half_adder ha6_35_2 (
.a(c5_34_2),.b(c5_34_1),.p(s6_35_2),.g(c6_35_2)
);
wire c6_36_1, s6_36_1;
full_adder fa6_36_1 (
.a(c4_35_1),.b(s5_36_2),.c(s5_36_1),.s(s6_36_1),.co(c6_36_1)
);
wire c6_36_2, s6_36_2;
half_adder ha6_36_2 (
.a(c5_35_2),.b(c5_35_1),.p(s6_36_2),.g(c6_36_2)
);
wire c6_37_1, s6_37_1;
full_adder fa6_37_1 (
.a(s5_37_2),.b(s5_37_1),.c(c5_36_2),.s(s6_37_1),.co(c6_37_1)
);
wire c6_38_1, s6_38_1;
full_adder fa6_38_1 (
.a(s5_38_2),.b(s5_38_1),.c(c5_37_2),.s(s6_38_1),.co(c6_38_1)
);
wire c6_39_1, s6_39_1;
full_adder fa6_39_1 (
.a(s5_39_2),.b(s5_39_1),.c(c5_38_2),.s(s6_39_1),.co(c6_39_1)
);
wire c6_40_1, s6_40_1;
full_adder fa6_40_1 (
.a(s5_40_2),.b(s5_40_1),.c(c5_39_2),.s(s6_40_1),.co(c6_40_1)
);
wire c6_41_1, s6_41_1;
full_adder fa6_41_1 (
.a(s5_41_2),.b(s5_41_1),.c(c5_40_2),.s(s6_41_1),.co(c6_41_1)
);
wire c6_42_1, s6_42_1;
full_adder fa6_42_1 (
.a(s5_42_2),.b(s5_42_1),.c(c5_41_2),.s(s6_42_1),.co(c6_42_1)
);
wire c6_43_1, s6_43_1;
full_adder fa6_43_1 (
.a(s5_43_2),.b(s5_43_1),.c(c5_42_2),.s(s6_43_1),.co(c6_43_1)
);
wire c6_44_1, s6_44_1;
full_adder fa6_44_1 (
.a(s5_44_2),.b(s5_44_1),.c(c5_43_2),.s(s6_44_1),.co(c6_44_1)
);
wire c6_45_1, s6_45_1;
full_adder fa6_45_1 (
.a(c4_44_1),.b(s5_45_1),.c(c5_44_2),.s(s6_45_1),.co(c6_45_1)
);
wire c6_46_1, s6_46_1;
full_adder fa6_46_1 (
.a(c4_45_1),.b(s5_46_1),.c(c5_45_1),.s(s6_46_1),.co(c6_46_1)
);
wire c6_47_1, s6_47_1;
full_adder fa6_47_1 (
.a(c4_46_1),.b(s5_47_1),.c(c5_46_1),.s(s6_47_1),.co(c6_47_1)
);
wire c6_48_1, s6_48_1;
full_adder fa6_48_1 (
.a(c4_47_1),.b(s5_48_1),.c(c5_47_1),.s(s6_48_1),.co(c6_48_1)
);
wire c6_49_1, s6_49_1;
full_adder fa6_49_1 (
.a(c4_48_1),.b(s5_49_1),.c(c5_48_1),.s(s6_49_1),.co(c6_49_1)
);
wire c6_50_1, s6_50_1;
full_adder fa6_50_1 (
.a(c4_49_1),.b(s5_50_1),.c(c5_49_1),.s(s6_50_1),.co(c6_50_1)
);
wire c6_51_1, s6_51_1;
full_adder fa6_51_1 (
.a(c4_50_1),.b(s5_51_1),.c(c5_50_1),.s(s6_51_1),.co(c6_51_1)
);
wire c6_52_1, s6_52_1;
half_adder ha6_52_1 (
.a(s5_52_1),.b(c5_51_1),.p(s6_52_1),.g(c6_52_1)
);
wire c6_53_1, s6_53_1;
half_adder ha6_53_1 (
.a(s5_53_1),.b(c5_52_1),.p(s6_53_1),.g(c6_53_1)
);
wire c6_54_1, s6_54_1;
half_adder ha6_54_1 (
.a(s5_54_1),.b(c5_53_1),.p(s6_54_1),.g(c6_54_1)
);
wire c6_55_1, s6_55_1;
half_adder ha6_55_1 (
.a(s5_55_1),.b(c5_54_1),.p(s6_55_1),.g(c6_55_1)
);
wire c6_56_1, s6_56_1;
half_adder ha6_56_1 (
.a(s5_56_1),.b(c5_55_1),.p(s6_56_1),.g(c6_56_1)
);
wire c6_57_1, s6_57_1;
half_adder ha6_57_1 (
.a(s5_57_1),.b(c5_56_1),.p(s6_57_1),.g(c6_57_1)
);
wire c6_58_1, s6_58_1;
half_adder ha6_58_1 (
.a(s5_58_1),.b(c5_57_1),.p(s6_58_1),.g(c6_58_1)
);
wire c6_59_1, s6_59_1;
half_adder ha6_59_1 (
.a(s5_59_1),.b(c5_58_1),.p(s6_59_1),.g(c6_59_1)
);
wire c6_60_1, s6_60_1;
half_adder ha6_60_1 (
.a(s5_60_1),.b(c5_59_1),.p(s6_60_1),.g(c6_60_1)
);
wire c6_61_1, s6_61_1;
half_adder ha6_61_1 (
.a(s5_61_1),.b(c5_60_1),.p(s6_61_1),.g(c6_61_1)
);
wire c6_62_1, s6_62_1;
half_adder ha6_62_1 (
.a(s5_62_1),.b(c5_61_1),.p(s6_62_1),.g(c6_62_1)
);
wire c6_63_1, s6_63_1;
half_adder ha6_63_1 (
.a(s5_63_1),.b(c5_62_1),.p(s6_63_1),.g(c6_63_1)
);
wire c7_7_1, s7_7_1;
half_adder ha7_7_1 (
.a(s6_7_1),.b(c6_6_1),.p(s7_7_1),.g(c7_7_1)
);
wire c7_8_1, s7_8_1;
half_adder ha7_8_1 (
.a(s6_8_1),.b(c6_7_1),.p(s7_8_1),.g(c7_8_1)
);
wire c7_9_1, s7_9_1;
half_adder ha7_9_1 (
.a(s6_9_1),.b(c6_8_1),.p(s7_9_1),.g(c7_9_1)
);
wire c7_10_1, s7_10_1;
half_adder ha7_10_1 (
.a(s6_10_1),.b(c6_9_1),.p(s7_10_1),.g(c7_10_1)
);
wire c7_11_1, s7_11_1;
half_adder ha7_11_1 (
.a(s6_11_1),.b(c6_10_1),.p(s7_11_1),.g(c7_11_1)
);
wire c7_12_1, s7_12_1;
half_adder ha7_12_1 (
.a(s6_12_1),.b(c6_11_1),.p(s7_12_1),.g(c7_12_1)
);
wire c7_13_1, s7_13_1;
half_adder ha7_13_1 (
.a(s6_13_1),.b(c6_12_1),.p(s7_13_1),.g(c7_13_1)
);
wire c7_14_1, s7_14_1;
half_adder ha7_14_1 (
.a(s6_14_1),.b(c6_13_1),.p(s7_14_1),.g(c7_14_1)
);
wire c7_15_1, s7_15_1;
half_adder ha7_15_1 (
.a(s6_15_1),.b(c6_14_1),.p(s7_15_1),.g(c7_15_1)
);
wire c7_16_1, s7_16_1;
half_adder ha7_16_1 (
.a(s6_16_1),.b(c6_15_1),.p(s7_16_1),.g(c7_16_1)
);
wire c7_17_1, s7_17_1;
half_adder ha7_17_1 (
.a(s6_17_1),.b(c6_16_1),.p(s7_17_1),.g(c7_17_1)
);
wire c7_18_1, s7_18_1;
half_adder ha7_18_1 (
.a(s6_18_1),.b(c6_17_1),.p(s7_18_1),.g(c7_18_1)
);
wire c7_19_1, s7_19_1;
half_adder ha7_19_1 (
.a(s6_19_1),.b(c6_18_1),.p(s7_19_1),.g(c7_19_1)
);
wire c7_20_1, s7_20_1;
half_adder ha7_20_1 (
.a(s6_20_1),.b(c6_19_1),.p(s7_20_1),.g(c7_20_1)
);
wire c7_21_1, s7_21_1;
half_adder ha7_21_1 (
.a(s6_21_1),.b(c6_20_1),.p(s7_21_1),.g(c7_21_1)
);
wire c7_22_1, s7_22_1;
full_adder fa7_22_1 (
.a(c5_21_1),.b(s6_22_1),.c(c6_21_1),.s(s7_22_1),.co(c7_22_1)
);
wire c7_23_1, s7_23_1;
full_adder fa7_23_1 (
.a(c5_22_1),.b(s6_23_1),.c(c6_22_1),.s(s7_23_1),.co(c7_23_1)
);
wire c7_24_1, s7_24_1;
full_adder fa7_24_1 (
.a(c5_23_1),.b(s6_24_1),.c(c6_23_1),.s(s7_24_1),.co(c7_24_1)
);
wire c7_25_1, s7_25_1;
full_adder fa7_25_1 (
.a(c5_24_1),.b(s6_25_1),.c(c6_24_1),.s(s7_25_1),.co(c7_25_1)
);
wire c7_26_1, s7_26_1;
full_adder fa7_26_1 (
.a(c5_25_1),.b(s6_26_1),.c(c6_25_1),.s(s7_26_1),.co(c7_26_1)
);
wire c7_27_1, s7_27_1;
full_adder fa7_27_1 (
.a(c5_26_1),.b(s6_27_1),.c(c6_26_1),.s(s7_27_1),.co(c7_27_1)
);
wire c7_28_1, s7_28_1;
full_adder fa7_28_1 (
.a(c5_27_1),.b(s6_28_1),.c(c6_27_1),.s(s7_28_1),.co(c7_28_1)
);
wire c7_29_1, s7_29_1;
full_adder fa7_29_1 (
.a(c5_28_1),.b(s6_29_1),.c(c6_28_1),.s(s7_29_1),.co(c7_29_1)
);
wire c7_30_1, s7_30_1;
full_adder fa7_30_1 (
.a(c5_29_1),.b(s6_30_1),.c(c6_29_1),.s(s7_30_1),.co(c7_30_1)
);
wire c7_31_1, s7_31_1;
full_adder fa7_31_1 (
.a(s6_31_2),.b(s6_31_1),.c(c6_30_1),.s(s7_31_1),.co(c7_31_1)
);
wire c7_32_1, s7_32_1;
full_adder fa7_32_1 (
.a(s6_32_2),.b(s6_32_1),.c(c6_31_2),.s(s7_32_1),.co(c7_32_1)
);
wire c7_33_1, s7_33_1;
full_adder fa7_33_1 (
.a(s6_33_2),.b(s6_33_1),.c(c6_32_2),.s(s7_33_1),.co(c7_33_1)
);
wire c7_34_1, s7_34_1;
full_adder fa7_34_1 (
.a(s6_34_2),.b(s6_34_1),.c(c6_33_2),.s(s7_34_1),.co(c7_34_1)
);
wire c7_35_1, s7_35_1;
full_adder fa7_35_1 (
.a(s6_35_2),.b(s6_35_1),.c(c6_34_2),.s(s7_35_1),.co(c7_35_1)
);
wire c7_36_1, s7_36_1;
full_adder fa7_36_1 (
.a(s6_36_2),.b(s6_36_1),.c(c6_35_2),.s(s7_36_1),.co(c7_36_1)
);
wire c7_37_1, s7_37_1;
full_adder fa7_37_1 (
.a(c5_36_1),.b(s6_37_1),.c(c6_36_2),.s(s7_37_1),.co(c7_37_1)
);
wire c7_38_1, s7_38_1;
full_adder fa7_38_1 (
.a(c5_37_1),.b(s6_38_1),.c(c6_37_1),.s(s7_38_1),.co(c7_38_1)
);
wire c7_39_1, s7_39_1;
full_adder fa7_39_1 (
.a(c5_38_1),.b(s6_39_1),.c(c6_38_1),.s(s7_39_1),.co(c7_39_1)
);
wire c7_40_1, s7_40_1;
full_adder fa7_40_1 (
.a(c5_39_1),.b(s6_40_1),.c(c6_39_1),.s(s7_40_1),.co(c7_40_1)
);
wire c7_41_1, s7_41_1;
full_adder fa7_41_1 (
.a(c5_40_1),.b(s6_41_1),.c(c6_40_1),.s(s7_41_1),.co(c7_41_1)
);
wire c7_42_1, s7_42_1;
full_adder fa7_42_1 (
.a(c5_41_1),.b(s6_42_1),.c(c6_41_1),.s(s7_42_1),.co(c7_42_1)
);
wire c7_43_1, s7_43_1;
full_adder fa7_43_1 (
.a(c5_42_1),.b(s6_43_1),.c(c6_42_1),.s(s7_43_1),.co(c7_43_1)
);
wire c7_44_1, s7_44_1;
full_adder fa7_44_1 (
.a(c5_43_1),.b(s6_44_1),.c(c6_43_1),.s(s7_44_1),.co(c7_44_1)
);
wire c7_45_1, s7_45_1;
full_adder fa7_45_1 (
.a(c5_44_1),.b(s6_45_1),.c(c6_44_1),.s(s7_45_1),.co(c7_45_1)
);
wire c7_46_1, s7_46_1;
half_adder ha7_46_1 (
.a(s6_46_1),.b(c6_45_1),.p(s7_46_1),.g(c7_46_1)
);
wire c7_47_1, s7_47_1;
half_adder ha7_47_1 (
.a(s6_47_1),.b(c6_46_1),.p(s7_47_1),.g(c7_47_1)
);
wire c7_48_1, s7_48_1;
half_adder ha7_48_1 (
.a(s6_48_1),.b(c6_47_1),.p(s7_48_1),.g(c7_48_1)
);
wire c7_49_1, s7_49_1;
half_adder ha7_49_1 (
.a(s6_49_1),.b(c6_48_1),.p(s7_49_1),.g(c7_49_1)
);
wire c7_50_1, s7_50_1;
half_adder ha7_50_1 (
.a(s6_50_1),.b(c6_49_1),.p(s7_50_1),.g(c7_50_1)
);
wire c7_51_1, s7_51_1;
half_adder ha7_51_1 (
.a(s6_51_1),.b(c6_50_1),.p(s7_51_1),.g(c7_51_1)
);
wire c7_52_1, s7_52_1;
half_adder ha7_52_1 (
.a(s6_52_1),.b(c6_51_1),.p(s7_52_1),.g(c7_52_1)
);
wire c7_53_1, s7_53_1;
half_adder ha7_53_1 (
.a(s6_53_1),.b(c6_52_1),.p(s7_53_1),.g(c7_53_1)
);
wire c7_54_1, s7_54_1;
half_adder ha7_54_1 (
.a(s6_54_1),.b(c6_53_1),.p(s7_54_1),.g(c7_54_1)
);
wire c7_55_1, s7_55_1;
half_adder ha7_55_1 (
.a(s6_55_1),.b(c6_54_1),.p(s7_55_1),.g(c7_55_1)
);
wire c7_56_1, s7_56_1;
half_adder ha7_56_1 (
.a(s6_56_1),.b(c6_55_1),.p(s7_56_1),.g(c7_56_1)
);
wire c7_57_1, s7_57_1;
half_adder ha7_57_1 (
.a(s6_57_1),.b(c6_56_1),.p(s7_57_1),.g(c7_57_1)
);
wire c7_58_1, s7_58_1;
half_adder ha7_58_1 (
.a(s6_58_1),.b(c6_57_1),.p(s7_58_1),.g(c7_58_1)
);
wire c7_59_1, s7_59_1;
half_adder ha7_59_1 (
.a(s6_59_1),.b(c6_58_1),.p(s7_59_1),.g(c7_59_1)
);
wire c7_60_1, s7_60_1;
half_adder ha7_60_1 (
.a(s6_60_1),.b(c6_59_1),.p(s7_60_1),.g(c7_60_1)
);
wire c7_61_1, s7_61_1;
half_adder ha7_61_1 (
.a(s6_61_1),.b(c6_60_1),.p(s7_61_1),.g(c7_61_1)
);
wire c7_62_1, s7_62_1;
half_adder ha7_62_1 (
.a(s6_62_1),.b(c6_61_1),.p(s7_62_1),.g(c7_62_1)
);
wire c7_63_1, s7_63_1;
half_adder ha7_63_1 (
.a(s6_63_1),.b(c6_62_1),.p(s7_63_1),.g(c7_63_1)
);
wire c8_8_1, s8_8_1;
half_adder ha8_8_1 (
.a(s7_8_1),.b(c7_7_1),.p(s8_8_1),.g(c8_8_1)
);
wire c8_9_1, s8_9_1;
half_adder ha8_9_1 (
.a(s7_9_1),.b(c7_8_1),.p(s8_9_1),.g(c8_9_1)
);
wire c8_10_1, s8_10_1;
half_adder ha8_10_1 (
.a(s7_10_1),.b(c7_9_1),.p(s8_10_1),.g(c8_10_1)
);
wire c8_11_1, s8_11_1;
half_adder ha8_11_1 (
.a(s7_11_1),.b(c7_10_1),.p(s8_11_1),.g(c8_11_1)
);
wire c8_12_1, s8_12_1;
half_adder ha8_12_1 (
.a(s7_12_1),.b(c7_11_1),.p(s8_12_1),.g(c8_12_1)
);
wire c8_13_1, s8_13_1;
half_adder ha8_13_1 (
.a(s7_13_1),.b(c7_12_1),.p(s8_13_1),.g(c8_13_1)
);
wire c8_14_1, s8_14_1;
half_adder ha8_14_1 (
.a(s7_14_1),.b(c7_13_1),.p(s8_14_1),.g(c8_14_1)
);
wire c8_15_1, s8_15_1;
half_adder ha8_15_1 (
.a(s7_15_1),.b(c7_14_1),.p(s8_15_1),.g(c8_15_1)
);
wire c8_16_1, s8_16_1;
half_adder ha8_16_1 (
.a(s7_16_1),.b(c7_15_1),.p(s8_16_1),.g(c8_16_1)
);
wire c8_17_1, s8_17_1;
half_adder ha8_17_1 (
.a(s7_17_1),.b(c7_16_1),.p(s8_17_1),.g(c8_17_1)
);
wire c8_18_1, s8_18_1;
half_adder ha8_18_1 (
.a(s7_18_1),.b(c7_17_1),.p(s8_18_1),.g(c8_18_1)
);
wire c8_19_1, s8_19_1;
half_adder ha8_19_1 (
.a(s7_19_1),.b(c7_18_1),.p(s8_19_1),.g(c8_19_1)
);
wire c8_20_1, s8_20_1;
half_adder ha8_20_1 (
.a(s7_20_1),.b(c7_19_1),.p(s8_20_1),.g(c8_20_1)
);
wire c8_21_1, s8_21_1;
half_adder ha8_21_1 (
.a(s7_21_1),.b(c7_20_1),.p(s8_21_1),.g(c8_21_1)
);
wire c8_22_1, s8_22_1;
half_adder ha8_22_1 (
.a(s7_22_1),.b(c7_21_1),.p(s8_22_1),.g(c8_22_1)
);
wire c8_23_1, s8_23_1;
half_adder ha8_23_1 (
.a(s7_23_1),.b(c7_22_1),.p(s8_23_1),.g(c8_23_1)
);
wire c8_24_1, s8_24_1;
half_adder ha8_24_1 (
.a(s7_24_1),.b(c7_23_1),.p(s8_24_1),.g(c8_24_1)
);
wire c8_25_1, s8_25_1;
half_adder ha8_25_1 (
.a(s7_25_1),.b(c7_24_1),.p(s8_25_1),.g(c8_25_1)
);
wire c8_26_1, s8_26_1;
half_adder ha8_26_1 (
.a(s7_26_1),.b(c7_25_1),.p(s8_26_1),.g(c8_26_1)
);
wire c8_27_1, s8_27_1;
half_adder ha8_27_1 (
.a(s7_27_1),.b(c7_26_1),.p(s8_27_1),.g(c8_27_1)
);
wire c8_28_1, s8_28_1;
half_adder ha8_28_1 (
.a(s7_28_1),.b(c7_27_1),.p(s8_28_1),.g(c8_28_1)
);
wire c8_29_1, s8_29_1;
half_adder ha8_29_1 (
.a(s7_29_1),.b(c7_28_1),.p(s8_29_1),.g(c8_29_1)
);
wire c8_30_1, s8_30_1;
half_adder ha8_30_1 (
.a(s7_30_1),.b(c7_29_1),.p(s8_30_1),.g(c8_30_1)
);
wire c8_31_1, s8_31_1;
half_adder ha8_31_1 (
.a(s7_31_1),.b(c7_30_1),.p(s8_31_1),.g(c8_31_1)
);
wire c8_32_1, s8_32_1;
full_adder fa8_32_1 (
.a(c6_31_1),.b(s7_32_1),.c(c7_31_1),.s(s8_32_1),.co(c8_32_1)
);
wire c8_33_1, s8_33_1;
full_adder fa8_33_1 (
.a(c6_32_1),.b(s7_33_1),.c(c7_32_1),.s(s8_33_1),.co(c8_33_1)
);
wire c8_34_1, s8_34_1;
full_adder fa8_34_1 (
.a(c6_33_1),.b(s7_34_1),.c(c7_33_1),.s(s8_34_1),.co(c8_34_1)
);
wire c8_35_1, s8_35_1;
full_adder fa8_35_1 (
.a(c6_34_1),.b(s7_35_1),.c(c7_34_1),.s(s8_35_1),.co(c8_35_1)
);
wire c8_36_1, s8_36_1;
full_adder fa8_36_1 (
.a(c6_35_1),.b(s7_36_1),.c(c7_35_1),.s(s8_36_1),.co(c8_36_1)
);
wire c8_37_1, s8_37_1;
full_adder fa8_37_1 (
.a(c6_36_1),.b(s7_37_1),.c(c7_36_1),.s(s8_37_1),.co(c8_37_1)
);
wire c8_38_1, s8_38_1;
half_adder ha8_38_1 (
.a(s7_38_1),.b(c7_37_1),.p(s8_38_1),.g(c8_38_1)
);
wire c8_39_1, s8_39_1;
half_adder ha8_39_1 (
.a(s7_39_1),.b(c7_38_1),.p(s8_39_1),.g(c8_39_1)
);
wire c8_40_1, s8_40_1;
half_adder ha8_40_1 (
.a(s7_40_1),.b(c7_39_1),.p(s8_40_1),.g(c8_40_1)
);
wire c8_41_1, s8_41_1;
half_adder ha8_41_1 (
.a(s7_41_1),.b(c7_40_1),.p(s8_41_1),.g(c8_41_1)
);
wire c8_42_1, s8_42_1;
half_adder ha8_42_1 (
.a(s7_42_1),.b(c7_41_1),.p(s8_42_1),.g(c8_42_1)
);
wire c8_43_1, s8_43_1;
half_adder ha8_43_1 (
.a(s7_43_1),.b(c7_42_1),.p(s8_43_1),.g(c8_43_1)
);
wire c8_44_1, s8_44_1;
half_adder ha8_44_1 (
.a(s7_44_1),.b(c7_43_1),.p(s8_44_1),.g(c8_44_1)
);
wire c8_45_1, s8_45_1;
half_adder ha8_45_1 (
.a(s7_45_1),.b(c7_44_1),.p(s8_45_1),.g(c8_45_1)
);
wire c8_46_1, s8_46_1;
half_adder ha8_46_1 (
.a(s7_46_1),.b(c7_45_1),.p(s8_46_1),.g(c8_46_1)
);
wire c8_47_1, s8_47_1;
half_adder ha8_47_1 (
.a(s7_47_1),.b(c7_46_1),.p(s8_47_1),.g(c8_47_1)
);
wire c8_48_1, s8_48_1;
half_adder ha8_48_1 (
.a(s7_48_1),.b(c7_47_1),.p(s8_48_1),.g(c8_48_1)
);
wire c8_49_1, s8_49_1;
half_adder ha8_49_1 (
.a(s7_49_1),.b(c7_48_1),.p(s8_49_1),.g(c8_49_1)
);
wire c8_50_1, s8_50_1;
half_adder ha8_50_1 (
.a(s7_50_1),.b(c7_49_1),.p(s8_50_1),.g(c8_50_1)
);
wire c8_51_1, s8_51_1;
half_adder ha8_51_1 (
.a(s7_51_1),.b(c7_50_1),.p(s8_51_1),.g(c8_51_1)
);
wire c8_52_1, s8_52_1;
half_adder ha8_52_1 (
.a(s7_52_1),.b(c7_51_1),.p(s8_52_1),.g(c8_52_1)
);
wire c8_53_1, s8_53_1;
half_adder ha8_53_1 (
.a(s7_53_1),.b(c7_52_1),.p(s8_53_1),.g(c8_53_1)
);
wire c8_54_1, s8_54_1;
half_adder ha8_54_1 (
.a(s7_54_1),.b(c7_53_1),.p(s8_54_1),.g(c8_54_1)
);
wire c8_55_1, s8_55_1;
half_adder ha8_55_1 (
.a(s7_55_1),.b(c7_54_1),.p(s8_55_1),.g(c8_55_1)
);
wire c8_56_1, s8_56_1;
half_adder ha8_56_1 (
.a(s7_56_1),.b(c7_55_1),.p(s8_56_1),.g(c8_56_1)
);
wire c8_57_1, s8_57_1;
half_adder ha8_57_1 (
.a(s7_57_1),.b(c7_56_1),.p(s8_57_1),.g(c8_57_1)
);
wire c8_58_1, s8_58_1;
half_adder ha8_58_1 (
.a(s7_58_1),.b(c7_57_1),.p(s8_58_1),.g(c8_58_1)
);
wire c8_59_1, s8_59_1;
half_adder ha8_59_1 (
.a(s7_59_1),.b(c7_58_1),.p(s8_59_1),.g(c8_59_1)
);
wire c8_60_1, s8_60_1;
half_adder ha8_60_1 (
.a(s7_60_1),.b(c7_59_1),.p(s8_60_1),.g(c8_60_1)
);
wire c8_61_1, s8_61_1;
half_adder ha8_61_1 (
.a(s7_61_1),.b(c7_60_1),.p(s8_61_1),.g(c8_61_1)
);
wire c8_62_1, s8_62_1;
half_adder ha8_62_1 (
.a(s7_62_1),.b(c7_61_1),.p(s8_62_1),.g(c8_62_1)
);
wire c8_63_1, s8_63_1;
half_adder ha8_63_1 (
.a(s7_63_1),.b(c7_62_1),.p(s8_63_1),.g(c8_63_1)
);
wire [63:0]A_t;
wire [63:0]B_t;
assign A_t[0] = 1'b0;
assign B_t[0] = A[0] & B[0];
assign A_t[1] = 1'b0;
assign B_t[1] = s1_1_1;
assign A_t[2] = 1'b0;
assign B_t[2] = s2_2_1;
assign A_t[3] = 1'b0;
assign B_t[3] = s3_3_1;
assign A_t[4] = 1'b0;
assign B_t[4] = s4_4_1;
assign A_t[5] = 1'b0;
assign B_t[5] = s5_5_1;
assign A_t[6] = 1'b0;
assign B_t[6] = s6_6_1;
assign A_t[7] = 1'b0;
assign B_t[7] = s7_7_1;
assign A_t[8] = 1'b0;
assign B_t[8] = s8_8_1;
assign A_t[9] = s8_9_1;
assign B_t[9] = c8_8_1;
assign A_t[10] = s8_10_1;
assign B_t[10] = c8_9_1;
assign A_t[11] = s8_11_1;
assign B_t[11] = c8_10_1;
assign A_t[12] = s8_12_1;
assign B_t[12] = c8_11_1;
assign A_t[13] = s8_13_1;
assign B_t[13] = c8_12_1;
assign A_t[14] = s8_14_1;
assign B_t[14] = c8_13_1;
assign A_t[15] = s8_15_1;
assign B_t[15] = c8_14_1;
assign A_t[16] = s8_16_1;
assign B_t[16] = c8_15_1;
assign A_t[17] = s8_17_1;
assign B_t[17] = c8_16_1;
assign A_t[18] = s8_18_1;
assign B_t[18] = c8_17_1;
assign A_t[19] = s8_19_1;
assign B_t[19] = c8_18_1;
assign A_t[20] = s8_20_1;
assign B_t[20] = c8_19_1;
assign A_t[21] = s8_21_1;
assign B_t[21] = c8_20_1;
assign A_t[22] = s8_22_1;
assign B_t[22] = c8_21_1;
assign A_t[23] = s8_23_1;
assign B_t[23] = c8_22_1;
assign A_t[24] = s8_24_1;
assign B_t[24] = c8_23_1;
assign A_t[25] = s8_25_1;
assign B_t[25] = c8_24_1;
assign A_t[26] = s8_26_1;
assign B_t[26] = c8_25_1;
assign A_t[27] = s8_27_1;
assign B_t[27] = c8_26_1;
assign A_t[28] = s8_28_1;
assign B_t[28] = c8_27_1;
assign A_t[29] = s8_29_1;
assign B_t[29] = c8_28_1;
assign A_t[30] = s8_30_1;
assign B_t[30] = c8_29_1;
assign A_t[31] = s8_31_1;
assign B_t[31] = c8_30_1;
assign A_t[32] = s8_32_1;
assign B_t[32] = c8_31_1;
assign A_t[33] = s8_33_1;
assign B_t[33] = c8_32_1;
assign A_t[34] = s8_34_1;
assign B_t[34] = c8_33_1;
assign A_t[35] = s8_35_1;
assign B_t[35] = c8_34_1;
assign A_t[36] = s8_36_1;
assign B_t[36] = c8_35_1;
assign A_t[37] = s8_37_1;
assign B_t[37] = c8_36_1;
assign A_t[38] = s8_38_1;
assign B_t[38] = c8_37_1;
assign A_t[39] = s8_39_1;
assign B_t[39] = c8_38_1;
assign A_t[40] = s8_40_1;
assign B_t[40] = c8_39_1;
assign A_t[41] = s8_41_1;
assign B_t[41] = c8_40_1;
assign A_t[42] = s8_42_1;
assign B_t[42] = c8_41_1;
assign A_t[43] = s8_43_1;
assign B_t[43] = c8_42_1;
assign A_t[44] = s8_44_1;
assign B_t[44] = c8_43_1;
assign A_t[45] = s8_45_1;
assign B_t[45] = c8_44_1;
assign A_t[46] = s8_46_1;
assign B_t[46] = c8_45_1;
assign A_t[47] = s8_47_1;
assign B_t[47] = c8_46_1;
assign A_t[48] = s8_48_1;
assign B_t[48] = c8_47_1;
assign A_t[49] = s8_49_1;
assign B_t[49] = c8_48_1;
assign A_t[50] = s8_50_1;
assign B_t[50] = c8_49_1;
assign A_t[51] = s8_51_1;
assign B_t[51] = c8_50_1;
assign A_t[52] = s8_52_1;
assign B_t[52] = c8_51_1;
assign A_t[53] = s8_53_1;
assign B_t[53] = c8_52_1;
assign A_t[54] = s8_54_1;
assign B_t[54] = c8_53_1;
assign A_t[55] = s8_55_1;
assign B_t[55] = c8_54_1;
assign A_t[56] = s8_56_1;
assign B_t[56] = c8_55_1;
assign A_t[57] = s8_57_1;
assign B_t[57] = c8_56_1;
assign A_t[58] = s8_58_1;
assign B_t[58] = c8_57_1;
assign A_t[59] = s8_59_1;
assign B_t[59] = c8_58_1;
assign A_t[60] = s8_60_1;
assign B_t[60] = c8_59_1;
assign A_t[61] = s8_61_1;
assign B_t[61] = c8_60_1;
assign A_t[62] = s8_62_1;
assign B_t[62] = c8_61_1;
assign A_t[63] = s8_63_1;
assign B_t[63] = c8_62_1;

adder64 Adder(
    .A(A_t), 
    .B(B_t), 
    .res(C), 
    .overflow()
    );

endmodule
