`define DEBUG